module Arbiter_1(
  input  [31:0] io_in_0_bits_data,
  output [31:0] io_out_bits_data
);
  assign io_out_bits_data = io_in_0_bits_data; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
