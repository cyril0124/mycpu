module Decoder(
  input  [31:0] io_inst,
  output        io_out_isBranch,
  output [1:0]  io_out_resultSrc,
  output        io_out_memWrEn,
  output [2:0]  io_out_memType,
  output [3:0]  io_out_aluOpSel,
  output        io_out_aluSrc,
  output [1:0]  io_out_immSrc,
  output        io_out_immSign,
  output        io_out_regWrEn
);
  wire [31:0] _decodeSigs_T = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_1 = 32'h3 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_3 = 32'h1003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_5 = 32'h2003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_7 = 32'h4003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_9 = 32'h5003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_11 = 32'h13 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [31:0] _decodeSigs_T_12 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_13 = 32'h1013 == _decodeSigs_T_12; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_15 = 32'h2013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_17 = 32'h3013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_19 = 32'h4013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_21 = 32'h5013 == _decodeSigs_T_12; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_23 = 32'h40005013 == _decodeSigs_T_12; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_25 = 32'h6013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_27 = 32'h7013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [31:0] _decodeSigs_T_28 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_29 = 32'h17 == _decodeSigs_T_28; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_31 = 32'h23 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_33 = 32'h1023 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_35 = 32'h2023 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [31:0] _decodeSigs_T_36 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_37 = 32'h33 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_39 = 32'h40000033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_41 = 32'h1033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_43 = 32'h2033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_45 = 32'h3033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_47 = 32'h4033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_49 = 32'h5033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_51 = 32'h40005033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_53 = 32'h6033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_55 = 32'h7033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_57 = 32'h37 == _decodeSigs_T_28; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_59 = 32'h63 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_61 = 32'h1063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_63 = 32'h4063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_65 = 32'h5063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_67 = 32'h6063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_69 = 32'h7063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_71 = 32'h67 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_73 = 32'h6f == _decodeSigs_T_28; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_75 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_77 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_88 = _decodeSigs_T_57 ? 1'h0 : _decodeSigs_T_59 | (_decodeSigs_T_61 | (_decodeSigs_T_63 | (
    _decodeSigs_T_65 | (_decodeSigs_T_67 | _decodeSigs_T_69)))); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_89 = _decodeSigs_T_55 ? 1'h0 : _decodeSigs_T_88; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_90 = _decodeSigs_T_53 ? 1'h0 : _decodeSigs_T_89; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_91 = _decodeSigs_T_51 ? 1'h0 : _decodeSigs_T_90; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_92 = _decodeSigs_T_49 ? 1'h0 : _decodeSigs_T_91; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_93 = _decodeSigs_T_47 ? 1'h0 : _decodeSigs_T_92; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_94 = _decodeSigs_T_45 ? 1'h0 : _decodeSigs_T_93; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_95 = _decodeSigs_T_43 ? 1'h0 : _decodeSigs_T_94; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_96 = _decodeSigs_T_41 ? 1'h0 : _decodeSigs_T_95; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_97 = _decodeSigs_T_39 ? 1'h0 : _decodeSigs_T_96; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_98 = _decodeSigs_T_37 ? 1'h0 : _decodeSigs_T_97; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_99 = _decodeSigs_T_35 ? 1'h0 : _decodeSigs_T_98; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_100 = _decodeSigs_T_33 ? 1'h0 : _decodeSigs_T_99; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_101 = _decodeSigs_T_31 ? 1'h0 : _decodeSigs_T_100; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_102 = _decodeSigs_T_29 ? 1'h0 : _decodeSigs_T_101; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_103 = _decodeSigs_T_27 ? 1'h0 : _decodeSigs_T_102; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_104 = _decodeSigs_T_25 ? 1'h0 : _decodeSigs_T_103; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_105 = _decodeSigs_T_23 ? 1'h0 : _decodeSigs_T_104; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_106 = _decodeSigs_T_21 ? 1'h0 : _decodeSigs_T_105; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_107 = _decodeSigs_T_19 ? 1'h0 : _decodeSigs_T_106; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_108 = _decodeSigs_T_17 ? 1'h0 : _decodeSigs_T_107; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_109 = _decodeSigs_T_15 ? 1'h0 : _decodeSigs_T_108; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_110 = _decodeSigs_T_13 ? 1'h0 : _decodeSigs_T_109; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_111 = _decodeSigs_T_11 ? 1'h0 : _decodeSigs_T_110; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_112 = _decodeSigs_T_9 ? 1'h0 : _decodeSigs_T_111; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_113 = _decodeSigs_T_7 ? 1'h0 : _decodeSigs_T_112; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_114 = _decodeSigs_T_5 ? 1'h0 : _decodeSigs_T_113; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_115 = _decodeSigs_T_3 ? 1'h0 : _decodeSigs_T_114; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_118 = _decodeSigs_T_73 ? 2'h2 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_119 = _decodeSigs_T_71 ? 2'h2 : _decodeSigs_T_118; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_120 = _decodeSigs_T_69 ? 2'h0 : _decodeSigs_T_119; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_121 = _decodeSigs_T_67 ? 2'h0 : _decodeSigs_T_120; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_122 = _decodeSigs_T_65 ? 2'h0 : _decodeSigs_T_121; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_123 = _decodeSigs_T_63 ? 2'h0 : _decodeSigs_T_122; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_124 = _decodeSigs_T_61 ? 2'h0 : _decodeSigs_T_123; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_125 = _decodeSigs_T_59 ? 2'h0 : _decodeSigs_T_124; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_126 = _decodeSigs_T_57 ? 2'h0 : _decodeSigs_T_125; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_127 = _decodeSigs_T_55 ? 2'h0 : _decodeSigs_T_126; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_128 = _decodeSigs_T_53 ? 2'h0 : _decodeSigs_T_127; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_129 = _decodeSigs_T_51 ? 2'h0 : _decodeSigs_T_128; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_130 = _decodeSigs_T_49 ? 2'h0 : _decodeSigs_T_129; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_131 = _decodeSigs_T_47 ? 2'h0 : _decodeSigs_T_130; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_132 = _decodeSigs_T_45 ? 2'h0 : _decodeSigs_T_131; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_133 = _decodeSigs_T_43 ? 2'h0 : _decodeSigs_T_132; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_134 = _decodeSigs_T_41 ? 2'h0 : _decodeSigs_T_133; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_135 = _decodeSigs_T_39 ? 2'h0 : _decodeSigs_T_134; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_136 = _decodeSigs_T_37 ? 2'h0 : _decodeSigs_T_135; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_137 = _decodeSigs_T_35 ? 2'h0 : _decodeSigs_T_136; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_138 = _decodeSigs_T_33 ? 2'h0 : _decodeSigs_T_137; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_139 = _decodeSigs_T_31 ? 2'h0 : _decodeSigs_T_138; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_140 = _decodeSigs_T_29 ? 2'h0 : _decodeSigs_T_139; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_141 = _decodeSigs_T_27 ? 2'h0 : _decodeSigs_T_140; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_142 = _decodeSigs_T_25 ? 2'h0 : _decodeSigs_T_141; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_143 = _decodeSigs_T_23 ? 2'h0 : _decodeSigs_T_142; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_144 = _decodeSigs_T_21 ? 2'h0 : _decodeSigs_T_143; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_145 = _decodeSigs_T_19 ? 2'h0 : _decodeSigs_T_144; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_146 = _decodeSigs_T_17 ? 2'h0 : _decodeSigs_T_145; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_147 = _decodeSigs_T_15 ? 2'h0 : _decodeSigs_T_146; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_148 = _decodeSigs_T_13 ? 2'h0 : _decodeSigs_T_147; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_149 = _decodeSigs_T_11 ? 2'h0 : _decodeSigs_T_148; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_150 = _decodeSigs_T_9 ? 2'h1 : _decodeSigs_T_149; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_151 = _decodeSigs_T_7 ? 2'h1 : _decodeSigs_T_150; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_152 = _decodeSigs_T_5 ? 2'h1 : _decodeSigs_T_151; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_153 = _decodeSigs_T_3 ? 2'h1 : _decodeSigs_T_152; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_178 = _decodeSigs_T_29 ? 1'h0 : _decodeSigs_T_31 | (_decodeSigs_T_33 | _decodeSigs_T_35); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_179 = _decodeSigs_T_27 ? 1'h0 : _decodeSigs_T_178; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_180 = _decodeSigs_T_25 ? 1'h0 : _decodeSigs_T_179; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_181 = _decodeSigs_T_23 ? 1'h0 : _decodeSigs_T_180; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_182 = _decodeSigs_T_21 ? 1'h0 : _decodeSigs_T_181; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_183 = _decodeSigs_T_19 ? 1'h0 : _decodeSigs_T_182; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_184 = _decodeSigs_T_17 ? 1'h0 : _decodeSigs_T_183; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_185 = _decodeSigs_T_15 ? 1'h0 : _decodeSigs_T_184; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_186 = _decodeSigs_T_13 ? 1'h0 : _decodeSigs_T_185; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_187 = _decodeSigs_T_11 ? 1'h0 : _decodeSigs_T_186; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_188 = _decodeSigs_T_9 ? 1'h0 : _decodeSigs_T_187; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_189 = _decodeSigs_T_7 ? 1'h0 : _decodeSigs_T_188; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_190 = _decodeSigs_T_5 ? 1'h0 : _decodeSigs_T_189; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_191 = _decodeSigs_T_3 ? 1'h0 : _decodeSigs_T_190; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_252 = _decodeSigs_T_33 ? 3'h1 : 3'h2; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_253 = _decodeSigs_T_31 ? 3'h0 : _decodeSigs_T_252; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_254 = _decodeSigs_T_29 ? 3'h2 : _decodeSigs_T_253; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_255 = _decodeSigs_T_27 ? 3'h2 : _decodeSigs_T_254; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_256 = _decodeSigs_T_25 ? 3'h2 : _decodeSigs_T_255; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_257 = _decodeSigs_T_23 ? 3'h2 : _decodeSigs_T_256; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_258 = _decodeSigs_T_21 ? 3'h2 : _decodeSigs_T_257; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_259 = _decodeSigs_T_19 ? 3'h2 : _decodeSigs_T_258; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_260 = _decodeSigs_T_17 ? 3'h2 : _decodeSigs_T_259; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_261 = _decodeSigs_T_15 ? 3'h2 : _decodeSigs_T_260; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_262 = _decodeSigs_T_13 ? 3'h2 : _decodeSigs_T_261; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_263 = _decodeSigs_T_11 ? 3'h2 : _decodeSigs_T_262; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_264 = _decodeSigs_T_9 ? 3'h1 : _decodeSigs_T_263; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_265 = _decodeSigs_T_7 ? 3'h0 : _decodeSigs_T_264; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_266 = _decodeSigs_T_5 ? 3'h2 : _decodeSigs_T_265; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_267 = _decodeSigs_T_3 ? 3'h1 : _decodeSigs_T_266; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_272 = _decodeSigs_T_69 ? 4'h7 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_273 = _decodeSigs_T_67 ? 4'h8 : _decodeSigs_T_272; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_274 = _decodeSigs_T_65 ? 4'h7 : _decodeSigs_T_273; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_275 = _decodeSigs_T_63 ? 4'h8 : _decodeSigs_T_274; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_276 = _decodeSigs_T_61 ? 4'h6 : _decodeSigs_T_275; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_277 = _decodeSigs_T_59 ? 4'h5 : _decodeSigs_T_276; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_278 = _decodeSigs_T_57 ? 4'he : _decodeSigs_T_277; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_279 = _decodeSigs_T_55 ? 4'h2 : _decodeSigs_T_278; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_280 = _decodeSigs_T_53 ? 4'h3 : _decodeSigs_T_279; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_281 = _decodeSigs_T_51 ? 4'hc : _decodeSigs_T_280; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_282 = _decodeSigs_T_49 ? 4'hb : _decodeSigs_T_281; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_283 = _decodeSigs_T_47 ? 4'h4 : _decodeSigs_T_282; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_284 = _decodeSigs_T_45 ? 4'h9 : _decodeSigs_T_283; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_285 = _decodeSigs_T_43 ? 4'h8 : _decodeSigs_T_284; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_286 = _decodeSigs_T_41 ? 4'ha : _decodeSigs_T_285; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_287 = _decodeSigs_T_39 ? 4'h1 : _decodeSigs_T_286; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_288 = _decodeSigs_T_37 ? 4'h0 : _decodeSigs_T_287; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_289 = _decodeSigs_T_35 ? 4'h0 : _decodeSigs_T_288; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_290 = _decodeSigs_T_33 ? 4'h0 : _decodeSigs_T_289; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_291 = _decodeSigs_T_31 ? 4'h0 : _decodeSigs_T_290; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_292 = _decodeSigs_T_29 ? 4'h0 : _decodeSigs_T_291; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_293 = _decodeSigs_T_27 ? 4'h2 : _decodeSigs_T_292; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_294 = _decodeSigs_T_25 ? 4'h3 : _decodeSigs_T_293; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_295 = _decodeSigs_T_23 ? 4'hc : _decodeSigs_T_294; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_296 = _decodeSigs_T_21 ? 4'hb : _decodeSigs_T_295; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_297 = _decodeSigs_T_19 ? 4'h4 : _decodeSigs_T_296; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_298 = _decodeSigs_T_17 ? 4'h9 : _decodeSigs_T_297; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_299 = _decodeSigs_T_15 ? 4'h8 : _decodeSigs_T_298; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_300 = _decodeSigs_T_13 ? 4'ha : _decodeSigs_T_299; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_301 = _decodeSigs_T_11 ? 4'h0 : _decodeSigs_T_300; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_302 = _decodeSigs_T_9 ? 4'h0 : _decodeSigs_T_301; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_303 = _decodeSigs_T_7 ? 4'h0 : _decodeSigs_T_302; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_304 = _decodeSigs_T_5 ? 4'h0 : _decodeSigs_T_303; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_305 = _decodeSigs_T_3 ? 4'h0 : _decodeSigs_T_304; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_310 = _decodeSigs_T_69 ? 1'h0 : _decodeSigs_T_71 | _decodeSigs_T_73; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_311 = _decodeSigs_T_67 ? 1'h0 : _decodeSigs_T_310; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_312 = _decodeSigs_T_65 ? 1'h0 : _decodeSigs_T_311; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_313 = _decodeSigs_T_63 ? 1'h0 : _decodeSigs_T_312; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_314 = _decodeSigs_T_61 ? 1'h0 : _decodeSigs_T_313; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_315 = _decodeSigs_T_59 ? 1'h0 : _decodeSigs_T_314; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_317 = _decodeSigs_T_55 ? 1'h0 : _decodeSigs_T_57 | _decodeSigs_T_315; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_318 = _decodeSigs_T_53 ? 1'h0 : _decodeSigs_T_317; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_319 = _decodeSigs_T_51 ? 1'h0 : _decodeSigs_T_318; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_320 = _decodeSigs_T_49 ? 1'h0 : _decodeSigs_T_319; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_321 = _decodeSigs_T_47 ? 1'h0 : _decodeSigs_T_320; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_322 = _decodeSigs_T_45 ? 1'h0 : _decodeSigs_T_321; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_323 = _decodeSigs_T_43 ? 1'h0 : _decodeSigs_T_322; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_324 = _decodeSigs_T_41 ? 1'h0 : _decodeSigs_T_323; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_325 = _decodeSigs_T_39 ? 1'h0 : _decodeSigs_T_324; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_326 = _decodeSigs_T_37 ? 1'h0 : _decodeSigs_T_325; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_346 = _decodeSigs_T_73 ? 3'h4 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_347 = _decodeSigs_T_71 ? 3'h0 : _decodeSigs_T_346; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_348 = _decodeSigs_T_69 ? 3'h2 : _decodeSigs_T_347; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_349 = _decodeSigs_T_67 ? 3'h2 : _decodeSigs_T_348; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_350 = _decodeSigs_T_65 ? 3'h2 : _decodeSigs_T_349; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_351 = _decodeSigs_T_63 ? 3'h2 : _decodeSigs_T_350; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_352 = _decodeSigs_T_61 ? 3'h2 : _decodeSigs_T_351; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_353 = _decodeSigs_T_59 ? 3'h2 : _decodeSigs_T_352; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_354 = _decodeSigs_T_57 ? 3'h3 : _decodeSigs_T_353; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_355 = _decodeSigs_T_55 ? 3'h0 : _decodeSigs_T_354; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_356 = _decodeSigs_T_53 ? 3'h0 : _decodeSigs_T_355; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_357 = _decodeSigs_T_51 ? 3'h0 : _decodeSigs_T_356; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_358 = _decodeSigs_T_49 ? 3'h0 : _decodeSigs_T_357; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_359 = _decodeSigs_T_47 ? 3'h0 : _decodeSigs_T_358; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_360 = _decodeSigs_T_45 ? 3'h0 : _decodeSigs_T_359; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_361 = _decodeSigs_T_43 ? 3'h0 : _decodeSigs_T_360; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_362 = _decodeSigs_T_41 ? 3'h0 : _decodeSigs_T_361; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_363 = _decodeSigs_T_39 ? 3'h0 : _decodeSigs_T_362; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_364 = _decodeSigs_T_37 ? 3'h0 : _decodeSigs_T_363; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_365 = _decodeSigs_T_35 ? 3'h1 : _decodeSigs_T_364; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_366 = _decodeSigs_T_33 ? 3'h1 : _decodeSigs_T_365; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_367 = _decodeSigs_T_31 ? 3'h1 : _decodeSigs_T_366; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_368 = _decodeSigs_T_29 ? 3'h3 : _decodeSigs_T_367; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_369 = _decodeSigs_T_27 ? 3'h0 : _decodeSigs_T_368; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_370 = _decodeSigs_T_25 ? 3'h0 : _decodeSigs_T_369; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_371 = _decodeSigs_T_23 ? 3'h0 : _decodeSigs_T_370; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_372 = _decodeSigs_T_21 ? 3'h0 : _decodeSigs_T_371; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_373 = _decodeSigs_T_19 ? 3'h0 : _decodeSigs_T_372; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_374 = _decodeSigs_T_17 ? 3'h0 : _decodeSigs_T_373; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_375 = _decodeSigs_T_15 ? 3'h0 : _decodeSigs_T_374; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_376 = _decodeSigs_T_13 ? 3'h0 : _decodeSigs_T_375; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_377 = _decodeSigs_T_11 ? 3'h0 : _decodeSigs_T_376; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_378 = _decodeSigs_T_9 ? 3'h0 : _decodeSigs_T_377; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_379 = _decodeSigs_T_7 ? 3'h0 : _decodeSigs_T_378; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_380 = _decodeSigs_T_5 ? 3'h0 : _decodeSigs_T_379; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_381 = _decodeSigs_T_3 ? 3'h0 : _decodeSigs_T_380; // @[Lookup.scala 34:39]
  wire [2:0] decodeSigs_7 = _decodeSigs_T_1 ? 3'h0 : _decodeSigs_T_381; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_382 = _decodeSigs_T_77 ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_383 = _decodeSigs_T_75 ? 1'h0 : _decodeSigs_T_382; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_384 = _decodeSigs_T_73 ? 1'h0 : _decodeSigs_T_383; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_386 = _decodeSigs_T_69 ? 1'h0 : _decodeSigs_T_71 | _decodeSigs_T_384; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_387 = _decodeSigs_T_67 ? 1'h0 : _decodeSigs_T_386; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_390 = _decodeSigs_T_61 ? 1'h0 : _decodeSigs_T_63 | (_decodeSigs_T_65 | _decodeSigs_T_387); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_391 = _decodeSigs_T_59 ? 1'h0 : _decodeSigs_T_390; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_392 = _decodeSigs_T_57 ? 1'h0 : _decodeSigs_T_391; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_393 = _decodeSigs_T_55 ? 1'h0 : _decodeSigs_T_392; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_394 = _decodeSigs_T_53 ? 1'h0 : _decodeSigs_T_393; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_395 = _decodeSigs_T_51 ? 1'h0 : _decodeSigs_T_394; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_396 = _decodeSigs_T_49 ? 1'h0 : _decodeSigs_T_395; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_397 = _decodeSigs_T_47 ? 1'h0 : _decodeSigs_T_396; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_398 = _decodeSigs_T_45 ? 1'h0 : _decodeSigs_T_397; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_399 = _decodeSigs_T_43 ? 1'h0 : _decodeSigs_T_398; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_400 = _decodeSigs_T_41 ? 1'h0 : _decodeSigs_T_399; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_401 = _decodeSigs_T_39 ? 1'h0 : _decodeSigs_T_400; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_402 = _decodeSigs_T_37 ? 1'h0 : _decodeSigs_T_401; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_406 = _decodeSigs_T_29 ? 1'h0 : _decodeSigs_T_31 | (_decodeSigs_T_33 | (_decodeSigs_T_35 |
    _decodeSigs_T_402)); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_410 = _decodeSigs_T_21 ? 1'h0 : _decodeSigs_T_23 | (_decodeSigs_T_25 | (_decodeSigs_T_27 |
    _decodeSigs_T_406)); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_414 = _decodeSigs_T_13 ? 1'h0 : _decodeSigs_T_15 | (_decodeSigs_T_17 | (_decodeSigs_T_19 |
    _decodeSigs_T_410)); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_416 = _decodeSigs_T_9 ? 1'h0 : _decodeSigs_T_11 | _decodeSigs_T_414; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_417 = _decodeSigs_T_7 ? 1'h0 : _decodeSigs_T_416; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_418 = _decodeSigs_T_5 ? 1'h0 : _decodeSigs_T_417; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_419 = _decodeSigs_T_3 ? 1'h0 : _decodeSigs_T_418; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_441 = _decodeSigs_T_35 ? 1'h0 : _decodeSigs_T_37 | (_decodeSigs_T_39 | (_decodeSigs_T_41 | (
    _decodeSigs_T_43 | (_decodeSigs_T_45 | (_decodeSigs_T_47 | (_decodeSigs_T_49 | (_decodeSigs_T_51 | (_decodeSigs_T_53
     | (_decodeSigs_T_55 | (_decodeSigs_T_57 | _decodeSigs_T_315)))))))))); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_442 = _decodeSigs_T_33 ? 1'h0 : _decodeSigs_T_441; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_443 = _decodeSigs_T_31 ? 1'h0 : _decodeSigs_T_442; // @[Lookup.scala 34:39]
  assign io_out_isBranch = _decodeSigs_T_1 ? 1'h0 : _decodeSigs_T_115; // @[Lookup.scala 34:39]
  assign io_out_resultSrc = _decodeSigs_T_1 ? 2'h1 : _decodeSigs_T_153; // @[Lookup.scala 34:39]
  assign io_out_memWrEn = _decodeSigs_T_1 ? 1'h0 : _decodeSigs_T_191; // @[Lookup.scala 34:39]
  assign io_out_memType = _decodeSigs_T_1 ? 3'h0 : _decodeSigs_T_267; // @[Lookup.scala 34:39]
  assign io_out_aluOpSel = _decodeSigs_T_1 ? 4'h0 : _decodeSigs_T_305; // @[Lookup.scala 34:39]
  assign io_out_aluSrc = _decodeSigs_T_1 | (_decodeSigs_T_3 | (_decodeSigs_T_5 | (_decodeSigs_T_7 | (_decodeSigs_T_9 | (
    _decodeSigs_T_11 | (_decodeSigs_T_13 | (_decodeSigs_T_15 | (_decodeSigs_T_17 | (_decodeSigs_T_19 | (_decodeSigs_T_21
     | (_decodeSigs_T_23 | (_decodeSigs_T_25 | (_decodeSigs_T_27 | (_decodeSigs_T_29 | (_decodeSigs_T_31 | (
    _decodeSigs_T_33 | (_decodeSigs_T_35 | _decodeSigs_T_326))))))))))))))))); // @[Lookup.scala 34:39]
  assign io_out_immSrc = decodeSigs_7[1:0]; // @[Decoder.scala 131:19]
  assign io_out_immSign = _decodeSigs_T_1 ? 1'h0 : _decodeSigs_T_419; // @[Lookup.scala 34:39]
  assign io_out_regWrEn = _decodeSigs_T_1 | (_decodeSigs_T_3 | (_decodeSigs_T_5 | (_decodeSigs_T_7 | (_decodeSigs_T_9 |
    (_decodeSigs_T_11 | (_decodeSigs_T_13 | (_decodeSigs_T_15 | (_decodeSigs_T_17 | (_decodeSigs_T_19 | (
    _decodeSigs_T_21 | (_decodeSigs_T_23 | (_decodeSigs_T_25 | (_decodeSigs_T_27 | (_decodeSigs_T_29 | _decodeSigs_T_443
    )))))))))))))); // @[Lookup.scala 34:39]
endmodule
