module BankRam1P_1_33(
  input        clock,
  input        reset,
  input  [6:0] io_addr,
  input        io_rw,
  input  [3:0] io_wmask,
  output [3:0] io_rdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg  ram_0 [0:127]; // @[SRAM.scala 36:26]
  wire  ram_0_io_rdata_MPORT_en; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_io_rdata_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_0_io_rdata_MPORT_data; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_1_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_1_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_1_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_1_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_2_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_2_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_2_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_2_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_3_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_3_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_3_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_3_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_4_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_4_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_4_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_4_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_5_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_5_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_5_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_5_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_6_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_6_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_6_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_6_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_7_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_7_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_7_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_7_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_8_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_8_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_8_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_8_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_9_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_9_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_9_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_9_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_10_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_10_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_10_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_10_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_11_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_11_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_11_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_11_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_12_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_12_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_12_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_12_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_13_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_13_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_13_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_13_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_14_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_14_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_14_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_14_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_15_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_15_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_15_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_15_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_16_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_16_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_16_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_16_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_17_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_17_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_17_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_17_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_18_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_18_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_18_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_18_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_19_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_19_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_19_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_19_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_20_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_20_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_20_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_20_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_21_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_21_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_21_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_21_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_22_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_22_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_22_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_22_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_23_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_23_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_23_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_23_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_24_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_24_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_24_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_24_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_25_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_25_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_25_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_25_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_26_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_26_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_26_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_26_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_27_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_27_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_27_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_27_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_28_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_28_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_28_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_28_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_29_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_29_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_29_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_29_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_30_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_30_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_30_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_30_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_31_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_31_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_31_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_31_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_32_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_32_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_32_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_32_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_33_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_33_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_33_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_33_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_34_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_34_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_34_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_34_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_35_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_35_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_35_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_35_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_36_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_36_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_36_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_36_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_37_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_37_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_37_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_37_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_38_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_38_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_38_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_38_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_39_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_39_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_39_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_39_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_40_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_40_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_40_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_40_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_41_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_41_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_41_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_41_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_42_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_42_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_42_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_42_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_43_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_43_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_43_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_43_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_44_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_44_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_44_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_44_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_45_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_45_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_45_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_45_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_46_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_46_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_46_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_46_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_47_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_47_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_47_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_47_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_48_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_48_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_48_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_48_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_49_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_49_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_49_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_49_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_50_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_50_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_50_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_50_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_51_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_51_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_51_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_51_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_52_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_52_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_52_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_52_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_53_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_53_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_53_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_53_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_54_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_54_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_54_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_54_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_55_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_55_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_55_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_55_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_56_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_56_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_56_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_56_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_57_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_57_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_57_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_57_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_58_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_58_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_58_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_58_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_59_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_59_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_59_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_59_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_60_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_60_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_60_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_60_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_61_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_61_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_61_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_61_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_62_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_62_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_62_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_62_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_63_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_63_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_63_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_63_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_64_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_64_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_64_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_64_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_65_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_65_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_65_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_65_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_66_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_66_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_66_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_66_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_67_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_67_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_67_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_67_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_68_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_68_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_68_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_68_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_69_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_69_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_69_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_69_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_70_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_70_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_70_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_70_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_71_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_71_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_71_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_71_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_72_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_72_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_72_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_72_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_73_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_73_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_73_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_73_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_74_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_74_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_74_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_74_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_75_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_75_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_75_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_75_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_76_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_76_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_76_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_76_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_77_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_77_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_77_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_77_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_78_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_78_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_78_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_78_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_79_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_79_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_79_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_79_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_80_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_80_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_80_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_80_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_81_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_81_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_81_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_81_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_82_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_82_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_82_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_82_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_83_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_83_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_83_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_83_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_84_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_84_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_84_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_84_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_85_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_85_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_85_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_85_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_86_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_86_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_86_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_86_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_87_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_87_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_87_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_87_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_88_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_88_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_88_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_88_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_89_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_89_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_89_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_89_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_90_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_90_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_90_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_90_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_91_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_91_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_91_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_91_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_92_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_92_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_92_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_92_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_93_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_93_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_93_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_93_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_94_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_94_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_94_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_94_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_95_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_95_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_95_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_95_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_96_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_96_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_96_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_96_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_97_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_97_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_97_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_97_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_98_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_98_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_98_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_98_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_99_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_99_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_99_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_99_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_100_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_100_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_100_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_100_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_101_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_101_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_101_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_101_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_102_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_102_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_102_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_102_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_103_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_103_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_103_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_103_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_104_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_104_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_104_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_104_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_105_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_105_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_105_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_105_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_106_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_106_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_106_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_106_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_107_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_107_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_107_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_107_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_108_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_108_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_108_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_108_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_109_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_109_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_109_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_109_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_110_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_110_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_110_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_110_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_111_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_111_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_111_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_111_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_112_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_112_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_112_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_112_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_113_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_113_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_113_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_113_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_114_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_114_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_114_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_114_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_115_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_115_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_115_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_115_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_116_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_116_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_116_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_116_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_117_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_117_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_117_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_117_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_118_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_118_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_118_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_118_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_119_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_119_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_119_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_119_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_120_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_120_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_120_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_120_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_121_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_121_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_121_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_121_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_122_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_122_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_122_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_122_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_123_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_123_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_123_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_123_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_124_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_124_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_124_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_124_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_125_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_125_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_125_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_125_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_126_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_126_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_126_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_126_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_127_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_127_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_127_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_127_en; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_128_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_0_MPORT_128_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_128_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_128_en; // @[SRAM.scala 36:26]
  reg  ram_0_io_rdata_MPORT_en_pipe_0;
  reg [6:0] ram_0_io_rdata_MPORT_addr_pipe_0;
  reg  ram_1 [0:127]; // @[SRAM.scala 36:26]
  wire  ram_1_io_rdata_MPORT_en; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_io_rdata_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_1_io_rdata_MPORT_data; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_1_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_1_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_1_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_1_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_2_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_2_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_2_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_2_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_3_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_3_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_3_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_3_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_4_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_4_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_4_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_4_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_5_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_5_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_5_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_5_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_6_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_6_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_6_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_6_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_7_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_7_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_7_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_7_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_8_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_8_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_8_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_8_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_9_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_9_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_9_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_9_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_10_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_10_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_10_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_10_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_11_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_11_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_11_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_11_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_12_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_12_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_12_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_12_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_13_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_13_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_13_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_13_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_14_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_14_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_14_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_14_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_15_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_15_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_15_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_15_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_16_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_16_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_16_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_16_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_17_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_17_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_17_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_17_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_18_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_18_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_18_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_18_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_19_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_19_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_19_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_19_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_20_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_20_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_20_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_20_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_21_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_21_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_21_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_21_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_22_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_22_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_22_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_22_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_23_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_23_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_23_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_23_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_24_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_24_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_24_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_24_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_25_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_25_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_25_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_25_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_26_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_26_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_26_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_26_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_27_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_27_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_27_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_27_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_28_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_28_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_28_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_28_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_29_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_29_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_29_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_29_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_30_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_30_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_30_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_30_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_31_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_31_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_31_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_31_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_32_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_32_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_32_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_32_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_33_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_33_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_33_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_33_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_34_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_34_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_34_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_34_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_35_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_35_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_35_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_35_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_36_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_36_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_36_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_36_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_37_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_37_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_37_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_37_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_38_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_38_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_38_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_38_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_39_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_39_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_39_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_39_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_40_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_40_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_40_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_40_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_41_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_41_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_41_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_41_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_42_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_42_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_42_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_42_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_43_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_43_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_43_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_43_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_44_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_44_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_44_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_44_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_45_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_45_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_45_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_45_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_46_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_46_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_46_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_46_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_47_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_47_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_47_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_47_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_48_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_48_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_48_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_48_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_49_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_49_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_49_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_49_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_50_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_50_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_50_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_50_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_51_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_51_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_51_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_51_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_52_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_52_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_52_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_52_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_53_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_53_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_53_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_53_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_54_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_54_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_54_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_54_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_55_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_55_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_55_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_55_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_56_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_56_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_56_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_56_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_57_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_57_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_57_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_57_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_58_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_58_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_58_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_58_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_59_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_59_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_59_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_59_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_60_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_60_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_60_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_60_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_61_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_61_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_61_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_61_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_62_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_62_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_62_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_62_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_63_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_63_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_63_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_63_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_64_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_64_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_64_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_64_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_65_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_65_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_65_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_65_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_66_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_66_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_66_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_66_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_67_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_67_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_67_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_67_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_68_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_68_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_68_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_68_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_69_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_69_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_69_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_69_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_70_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_70_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_70_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_70_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_71_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_71_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_71_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_71_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_72_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_72_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_72_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_72_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_73_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_73_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_73_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_73_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_74_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_74_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_74_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_74_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_75_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_75_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_75_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_75_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_76_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_76_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_76_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_76_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_77_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_77_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_77_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_77_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_78_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_78_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_78_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_78_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_79_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_79_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_79_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_79_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_80_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_80_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_80_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_80_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_81_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_81_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_81_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_81_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_82_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_82_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_82_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_82_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_83_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_83_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_83_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_83_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_84_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_84_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_84_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_84_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_85_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_85_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_85_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_85_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_86_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_86_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_86_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_86_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_87_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_87_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_87_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_87_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_88_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_88_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_88_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_88_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_89_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_89_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_89_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_89_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_90_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_90_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_90_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_90_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_91_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_91_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_91_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_91_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_92_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_92_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_92_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_92_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_93_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_93_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_93_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_93_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_94_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_94_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_94_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_94_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_95_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_95_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_95_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_95_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_96_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_96_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_96_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_96_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_97_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_97_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_97_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_97_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_98_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_98_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_98_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_98_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_99_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_99_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_99_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_99_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_100_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_100_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_100_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_100_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_101_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_101_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_101_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_101_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_102_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_102_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_102_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_102_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_103_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_103_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_103_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_103_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_104_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_104_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_104_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_104_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_105_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_105_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_105_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_105_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_106_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_106_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_106_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_106_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_107_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_107_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_107_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_107_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_108_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_108_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_108_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_108_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_109_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_109_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_109_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_109_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_110_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_110_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_110_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_110_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_111_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_111_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_111_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_111_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_112_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_112_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_112_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_112_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_113_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_113_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_113_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_113_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_114_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_114_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_114_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_114_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_115_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_115_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_115_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_115_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_116_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_116_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_116_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_116_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_117_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_117_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_117_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_117_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_118_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_118_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_118_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_118_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_119_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_119_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_119_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_119_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_120_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_120_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_120_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_120_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_121_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_121_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_121_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_121_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_122_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_122_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_122_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_122_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_123_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_123_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_123_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_123_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_124_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_124_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_124_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_124_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_125_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_125_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_125_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_125_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_126_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_126_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_126_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_126_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_127_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_127_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_127_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_127_en; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_128_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_1_MPORT_128_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_128_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_128_en; // @[SRAM.scala 36:26]
  reg  ram_1_io_rdata_MPORT_en_pipe_0;
  reg [6:0] ram_1_io_rdata_MPORT_addr_pipe_0;
  reg  ram_2 [0:127]; // @[SRAM.scala 36:26]
  wire  ram_2_io_rdata_MPORT_en; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_io_rdata_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_2_io_rdata_MPORT_data; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_1_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_1_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_1_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_1_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_2_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_2_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_2_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_2_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_3_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_3_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_3_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_3_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_4_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_4_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_4_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_4_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_5_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_5_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_5_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_5_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_6_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_6_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_6_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_6_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_7_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_7_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_7_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_7_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_8_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_8_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_8_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_8_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_9_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_9_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_9_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_9_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_10_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_10_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_10_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_10_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_11_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_11_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_11_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_11_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_12_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_12_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_12_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_12_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_13_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_13_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_13_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_13_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_14_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_14_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_14_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_14_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_15_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_15_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_15_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_15_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_16_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_16_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_16_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_16_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_17_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_17_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_17_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_17_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_18_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_18_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_18_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_18_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_19_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_19_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_19_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_19_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_20_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_20_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_20_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_20_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_21_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_21_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_21_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_21_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_22_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_22_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_22_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_22_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_23_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_23_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_23_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_23_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_24_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_24_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_24_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_24_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_25_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_25_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_25_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_25_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_26_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_26_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_26_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_26_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_27_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_27_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_27_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_27_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_28_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_28_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_28_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_28_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_29_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_29_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_29_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_29_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_30_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_30_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_30_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_30_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_31_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_31_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_31_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_31_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_32_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_32_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_32_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_32_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_33_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_33_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_33_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_33_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_34_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_34_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_34_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_34_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_35_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_35_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_35_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_35_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_36_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_36_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_36_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_36_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_37_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_37_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_37_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_37_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_38_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_38_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_38_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_38_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_39_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_39_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_39_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_39_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_40_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_40_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_40_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_40_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_41_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_41_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_41_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_41_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_42_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_42_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_42_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_42_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_43_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_43_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_43_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_43_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_44_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_44_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_44_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_44_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_45_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_45_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_45_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_45_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_46_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_46_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_46_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_46_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_47_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_47_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_47_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_47_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_48_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_48_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_48_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_48_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_49_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_49_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_49_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_49_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_50_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_50_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_50_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_50_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_51_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_51_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_51_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_51_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_52_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_52_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_52_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_52_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_53_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_53_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_53_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_53_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_54_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_54_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_54_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_54_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_55_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_55_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_55_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_55_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_56_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_56_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_56_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_56_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_57_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_57_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_57_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_57_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_58_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_58_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_58_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_58_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_59_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_59_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_59_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_59_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_60_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_60_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_60_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_60_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_61_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_61_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_61_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_61_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_62_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_62_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_62_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_62_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_63_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_63_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_63_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_63_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_64_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_64_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_64_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_64_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_65_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_65_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_65_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_65_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_66_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_66_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_66_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_66_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_67_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_67_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_67_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_67_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_68_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_68_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_68_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_68_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_69_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_69_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_69_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_69_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_70_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_70_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_70_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_70_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_71_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_71_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_71_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_71_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_72_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_72_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_72_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_72_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_73_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_73_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_73_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_73_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_74_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_74_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_74_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_74_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_75_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_75_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_75_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_75_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_76_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_76_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_76_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_76_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_77_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_77_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_77_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_77_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_78_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_78_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_78_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_78_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_79_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_79_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_79_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_79_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_80_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_80_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_80_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_80_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_81_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_81_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_81_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_81_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_82_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_82_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_82_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_82_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_83_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_83_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_83_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_83_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_84_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_84_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_84_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_84_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_85_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_85_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_85_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_85_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_86_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_86_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_86_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_86_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_87_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_87_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_87_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_87_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_88_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_88_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_88_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_88_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_89_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_89_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_89_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_89_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_90_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_90_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_90_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_90_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_91_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_91_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_91_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_91_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_92_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_92_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_92_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_92_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_93_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_93_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_93_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_93_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_94_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_94_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_94_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_94_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_95_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_95_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_95_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_95_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_96_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_96_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_96_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_96_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_97_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_97_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_97_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_97_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_98_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_98_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_98_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_98_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_99_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_99_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_99_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_99_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_100_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_100_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_100_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_100_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_101_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_101_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_101_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_101_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_102_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_102_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_102_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_102_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_103_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_103_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_103_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_103_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_104_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_104_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_104_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_104_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_105_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_105_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_105_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_105_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_106_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_106_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_106_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_106_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_107_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_107_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_107_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_107_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_108_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_108_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_108_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_108_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_109_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_109_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_109_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_109_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_110_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_110_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_110_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_110_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_111_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_111_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_111_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_111_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_112_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_112_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_112_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_112_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_113_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_113_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_113_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_113_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_114_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_114_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_114_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_114_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_115_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_115_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_115_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_115_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_116_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_116_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_116_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_116_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_117_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_117_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_117_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_117_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_118_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_118_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_118_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_118_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_119_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_119_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_119_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_119_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_120_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_120_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_120_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_120_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_121_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_121_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_121_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_121_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_122_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_122_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_122_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_122_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_123_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_123_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_123_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_123_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_124_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_124_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_124_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_124_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_125_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_125_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_125_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_125_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_126_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_126_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_126_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_126_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_127_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_127_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_127_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_127_en; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_128_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_2_MPORT_128_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_128_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_128_en; // @[SRAM.scala 36:26]
  reg  ram_2_io_rdata_MPORT_en_pipe_0;
  reg [6:0] ram_2_io_rdata_MPORT_addr_pipe_0;
  reg  ram_3 [0:127]; // @[SRAM.scala 36:26]
  wire  ram_3_io_rdata_MPORT_en; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_io_rdata_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_3_io_rdata_MPORT_data; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_1_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_1_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_1_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_1_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_2_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_2_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_2_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_2_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_3_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_3_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_3_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_3_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_4_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_4_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_4_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_4_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_5_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_5_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_5_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_5_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_6_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_6_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_6_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_6_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_7_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_7_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_7_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_7_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_8_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_8_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_8_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_8_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_9_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_9_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_9_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_9_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_10_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_10_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_10_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_10_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_11_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_11_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_11_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_11_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_12_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_12_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_12_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_12_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_13_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_13_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_13_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_13_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_14_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_14_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_14_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_14_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_15_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_15_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_15_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_15_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_16_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_16_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_16_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_16_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_17_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_17_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_17_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_17_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_18_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_18_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_18_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_18_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_19_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_19_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_19_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_19_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_20_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_20_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_20_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_20_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_21_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_21_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_21_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_21_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_22_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_22_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_22_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_22_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_23_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_23_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_23_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_23_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_24_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_24_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_24_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_24_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_25_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_25_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_25_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_25_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_26_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_26_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_26_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_26_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_27_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_27_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_27_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_27_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_28_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_28_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_28_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_28_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_29_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_29_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_29_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_29_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_30_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_30_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_30_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_30_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_31_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_31_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_31_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_31_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_32_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_32_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_32_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_32_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_33_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_33_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_33_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_33_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_34_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_34_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_34_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_34_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_35_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_35_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_35_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_35_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_36_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_36_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_36_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_36_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_37_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_37_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_37_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_37_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_38_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_38_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_38_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_38_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_39_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_39_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_39_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_39_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_40_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_40_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_40_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_40_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_41_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_41_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_41_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_41_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_42_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_42_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_42_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_42_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_43_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_43_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_43_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_43_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_44_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_44_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_44_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_44_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_45_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_45_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_45_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_45_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_46_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_46_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_46_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_46_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_47_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_47_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_47_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_47_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_48_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_48_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_48_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_48_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_49_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_49_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_49_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_49_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_50_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_50_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_50_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_50_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_51_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_51_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_51_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_51_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_52_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_52_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_52_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_52_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_53_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_53_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_53_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_53_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_54_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_54_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_54_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_54_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_55_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_55_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_55_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_55_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_56_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_56_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_56_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_56_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_57_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_57_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_57_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_57_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_58_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_58_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_58_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_58_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_59_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_59_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_59_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_59_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_60_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_60_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_60_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_60_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_61_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_61_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_61_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_61_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_62_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_62_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_62_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_62_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_63_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_63_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_63_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_63_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_64_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_64_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_64_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_64_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_65_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_65_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_65_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_65_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_66_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_66_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_66_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_66_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_67_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_67_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_67_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_67_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_68_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_68_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_68_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_68_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_69_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_69_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_69_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_69_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_70_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_70_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_70_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_70_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_71_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_71_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_71_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_71_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_72_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_72_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_72_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_72_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_73_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_73_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_73_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_73_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_74_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_74_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_74_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_74_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_75_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_75_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_75_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_75_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_76_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_76_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_76_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_76_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_77_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_77_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_77_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_77_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_78_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_78_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_78_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_78_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_79_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_79_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_79_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_79_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_80_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_80_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_80_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_80_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_81_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_81_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_81_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_81_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_82_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_82_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_82_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_82_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_83_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_83_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_83_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_83_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_84_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_84_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_84_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_84_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_85_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_85_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_85_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_85_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_86_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_86_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_86_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_86_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_87_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_87_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_87_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_87_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_88_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_88_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_88_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_88_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_89_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_89_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_89_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_89_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_90_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_90_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_90_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_90_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_91_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_91_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_91_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_91_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_92_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_92_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_92_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_92_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_93_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_93_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_93_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_93_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_94_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_94_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_94_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_94_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_95_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_95_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_95_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_95_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_96_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_96_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_96_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_96_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_97_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_97_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_97_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_97_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_98_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_98_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_98_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_98_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_99_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_99_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_99_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_99_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_100_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_100_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_100_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_100_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_101_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_101_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_101_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_101_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_102_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_102_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_102_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_102_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_103_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_103_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_103_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_103_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_104_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_104_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_104_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_104_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_105_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_105_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_105_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_105_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_106_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_106_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_106_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_106_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_107_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_107_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_107_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_107_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_108_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_108_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_108_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_108_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_109_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_109_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_109_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_109_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_110_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_110_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_110_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_110_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_111_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_111_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_111_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_111_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_112_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_112_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_112_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_112_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_113_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_113_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_113_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_113_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_114_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_114_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_114_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_114_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_115_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_115_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_115_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_115_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_116_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_116_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_116_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_116_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_117_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_117_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_117_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_117_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_118_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_118_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_118_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_118_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_119_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_119_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_119_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_119_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_120_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_120_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_120_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_120_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_121_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_121_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_121_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_121_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_122_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_122_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_122_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_122_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_123_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_123_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_123_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_123_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_124_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_124_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_124_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_124_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_125_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_125_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_125_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_125_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_126_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_126_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_126_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_126_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_127_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_127_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_127_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_127_en; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_128_data; // @[SRAM.scala 36:26]
  wire [6:0] ram_3_MPORT_128_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_128_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_128_en; // @[SRAM.scala 36:26]
  reg  ram_3_io_rdata_MPORT_en_pipe_0;
  reg [6:0] ram_3_io_rdata_MPORT_addr_pipe_0;
  wire [1:0] io_rdata_lo = {ram_1_io_rdata_MPORT_data,ram_0_io_rdata_MPORT_data}; // @[SRAM.scala 75:39]
  wire [1:0] io_rdata_hi = {ram_3_io_rdata_MPORT_data,ram_2_io_rdata_MPORT_data}; // @[SRAM.scala 75:39]
  assign ram_0_io_rdata_MPORT_en = ram_0_io_rdata_MPORT_en_pipe_0;
  assign ram_0_io_rdata_MPORT_addr = ram_0_io_rdata_MPORT_addr_pipe_0;
  assign ram_0_io_rdata_MPORT_data = ram_0[ram_0_io_rdata_MPORT_addr]; // @[SRAM.scala 36:26]
  assign ram_0_MPORT_data = 1'h0;
  assign ram_0_MPORT_addr = 7'h0;
  assign ram_0_MPORT_mask = 1'h1;
  assign ram_0_MPORT_en = reset;
  assign ram_0_MPORT_1_data = 1'h0;
  assign ram_0_MPORT_1_addr = 7'h1;
  assign ram_0_MPORT_1_mask = 1'h1;
  assign ram_0_MPORT_1_en = reset;
  assign ram_0_MPORT_2_data = 1'h0;
  assign ram_0_MPORT_2_addr = 7'h2;
  assign ram_0_MPORT_2_mask = 1'h1;
  assign ram_0_MPORT_2_en = reset;
  assign ram_0_MPORT_3_data = 1'h0;
  assign ram_0_MPORT_3_addr = 7'h3;
  assign ram_0_MPORT_3_mask = 1'h1;
  assign ram_0_MPORT_3_en = reset;
  assign ram_0_MPORT_4_data = 1'h0;
  assign ram_0_MPORT_4_addr = 7'h4;
  assign ram_0_MPORT_4_mask = 1'h1;
  assign ram_0_MPORT_4_en = reset;
  assign ram_0_MPORT_5_data = 1'h0;
  assign ram_0_MPORT_5_addr = 7'h5;
  assign ram_0_MPORT_5_mask = 1'h1;
  assign ram_0_MPORT_5_en = reset;
  assign ram_0_MPORT_6_data = 1'h0;
  assign ram_0_MPORT_6_addr = 7'h6;
  assign ram_0_MPORT_6_mask = 1'h1;
  assign ram_0_MPORT_6_en = reset;
  assign ram_0_MPORT_7_data = 1'h0;
  assign ram_0_MPORT_7_addr = 7'h7;
  assign ram_0_MPORT_7_mask = 1'h1;
  assign ram_0_MPORT_7_en = reset;
  assign ram_0_MPORT_8_data = 1'h0;
  assign ram_0_MPORT_8_addr = 7'h8;
  assign ram_0_MPORT_8_mask = 1'h1;
  assign ram_0_MPORT_8_en = reset;
  assign ram_0_MPORT_9_data = 1'h0;
  assign ram_0_MPORT_9_addr = 7'h9;
  assign ram_0_MPORT_9_mask = 1'h1;
  assign ram_0_MPORT_9_en = reset;
  assign ram_0_MPORT_10_data = 1'h0;
  assign ram_0_MPORT_10_addr = 7'ha;
  assign ram_0_MPORT_10_mask = 1'h1;
  assign ram_0_MPORT_10_en = reset;
  assign ram_0_MPORT_11_data = 1'h0;
  assign ram_0_MPORT_11_addr = 7'hb;
  assign ram_0_MPORT_11_mask = 1'h1;
  assign ram_0_MPORT_11_en = reset;
  assign ram_0_MPORT_12_data = 1'h0;
  assign ram_0_MPORT_12_addr = 7'hc;
  assign ram_0_MPORT_12_mask = 1'h1;
  assign ram_0_MPORT_12_en = reset;
  assign ram_0_MPORT_13_data = 1'h0;
  assign ram_0_MPORT_13_addr = 7'hd;
  assign ram_0_MPORT_13_mask = 1'h1;
  assign ram_0_MPORT_13_en = reset;
  assign ram_0_MPORT_14_data = 1'h0;
  assign ram_0_MPORT_14_addr = 7'he;
  assign ram_0_MPORT_14_mask = 1'h1;
  assign ram_0_MPORT_14_en = reset;
  assign ram_0_MPORT_15_data = 1'h0;
  assign ram_0_MPORT_15_addr = 7'hf;
  assign ram_0_MPORT_15_mask = 1'h1;
  assign ram_0_MPORT_15_en = reset;
  assign ram_0_MPORT_16_data = 1'h0;
  assign ram_0_MPORT_16_addr = 7'h10;
  assign ram_0_MPORT_16_mask = 1'h1;
  assign ram_0_MPORT_16_en = reset;
  assign ram_0_MPORT_17_data = 1'h0;
  assign ram_0_MPORT_17_addr = 7'h11;
  assign ram_0_MPORT_17_mask = 1'h1;
  assign ram_0_MPORT_17_en = reset;
  assign ram_0_MPORT_18_data = 1'h0;
  assign ram_0_MPORT_18_addr = 7'h12;
  assign ram_0_MPORT_18_mask = 1'h1;
  assign ram_0_MPORT_18_en = reset;
  assign ram_0_MPORT_19_data = 1'h0;
  assign ram_0_MPORT_19_addr = 7'h13;
  assign ram_0_MPORT_19_mask = 1'h1;
  assign ram_0_MPORT_19_en = reset;
  assign ram_0_MPORT_20_data = 1'h0;
  assign ram_0_MPORT_20_addr = 7'h14;
  assign ram_0_MPORT_20_mask = 1'h1;
  assign ram_0_MPORT_20_en = reset;
  assign ram_0_MPORT_21_data = 1'h0;
  assign ram_0_MPORT_21_addr = 7'h15;
  assign ram_0_MPORT_21_mask = 1'h1;
  assign ram_0_MPORT_21_en = reset;
  assign ram_0_MPORT_22_data = 1'h0;
  assign ram_0_MPORT_22_addr = 7'h16;
  assign ram_0_MPORT_22_mask = 1'h1;
  assign ram_0_MPORT_22_en = reset;
  assign ram_0_MPORT_23_data = 1'h0;
  assign ram_0_MPORT_23_addr = 7'h17;
  assign ram_0_MPORT_23_mask = 1'h1;
  assign ram_0_MPORT_23_en = reset;
  assign ram_0_MPORT_24_data = 1'h0;
  assign ram_0_MPORT_24_addr = 7'h18;
  assign ram_0_MPORT_24_mask = 1'h1;
  assign ram_0_MPORT_24_en = reset;
  assign ram_0_MPORT_25_data = 1'h0;
  assign ram_0_MPORT_25_addr = 7'h19;
  assign ram_0_MPORT_25_mask = 1'h1;
  assign ram_0_MPORT_25_en = reset;
  assign ram_0_MPORT_26_data = 1'h0;
  assign ram_0_MPORT_26_addr = 7'h1a;
  assign ram_0_MPORT_26_mask = 1'h1;
  assign ram_0_MPORT_26_en = reset;
  assign ram_0_MPORT_27_data = 1'h0;
  assign ram_0_MPORT_27_addr = 7'h1b;
  assign ram_0_MPORT_27_mask = 1'h1;
  assign ram_0_MPORT_27_en = reset;
  assign ram_0_MPORT_28_data = 1'h0;
  assign ram_0_MPORT_28_addr = 7'h1c;
  assign ram_0_MPORT_28_mask = 1'h1;
  assign ram_0_MPORT_28_en = reset;
  assign ram_0_MPORT_29_data = 1'h0;
  assign ram_0_MPORT_29_addr = 7'h1d;
  assign ram_0_MPORT_29_mask = 1'h1;
  assign ram_0_MPORT_29_en = reset;
  assign ram_0_MPORT_30_data = 1'h0;
  assign ram_0_MPORT_30_addr = 7'h1e;
  assign ram_0_MPORT_30_mask = 1'h1;
  assign ram_0_MPORT_30_en = reset;
  assign ram_0_MPORT_31_data = 1'h0;
  assign ram_0_MPORT_31_addr = 7'h1f;
  assign ram_0_MPORT_31_mask = 1'h1;
  assign ram_0_MPORT_31_en = reset;
  assign ram_0_MPORT_32_data = 1'h0;
  assign ram_0_MPORT_32_addr = 7'h20;
  assign ram_0_MPORT_32_mask = 1'h1;
  assign ram_0_MPORT_32_en = reset;
  assign ram_0_MPORT_33_data = 1'h0;
  assign ram_0_MPORT_33_addr = 7'h21;
  assign ram_0_MPORT_33_mask = 1'h1;
  assign ram_0_MPORT_33_en = reset;
  assign ram_0_MPORT_34_data = 1'h0;
  assign ram_0_MPORT_34_addr = 7'h22;
  assign ram_0_MPORT_34_mask = 1'h1;
  assign ram_0_MPORT_34_en = reset;
  assign ram_0_MPORT_35_data = 1'h0;
  assign ram_0_MPORT_35_addr = 7'h23;
  assign ram_0_MPORT_35_mask = 1'h1;
  assign ram_0_MPORT_35_en = reset;
  assign ram_0_MPORT_36_data = 1'h0;
  assign ram_0_MPORT_36_addr = 7'h24;
  assign ram_0_MPORT_36_mask = 1'h1;
  assign ram_0_MPORT_36_en = reset;
  assign ram_0_MPORT_37_data = 1'h0;
  assign ram_0_MPORT_37_addr = 7'h25;
  assign ram_0_MPORT_37_mask = 1'h1;
  assign ram_0_MPORT_37_en = reset;
  assign ram_0_MPORT_38_data = 1'h0;
  assign ram_0_MPORT_38_addr = 7'h26;
  assign ram_0_MPORT_38_mask = 1'h1;
  assign ram_0_MPORT_38_en = reset;
  assign ram_0_MPORT_39_data = 1'h0;
  assign ram_0_MPORT_39_addr = 7'h27;
  assign ram_0_MPORT_39_mask = 1'h1;
  assign ram_0_MPORT_39_en = reset;
  assign ram_0_MPORT_40_data = 1'h0;
  assign ram_0_MPORT_40_addr = 7'h28;
  assign ram_0_MPORT_40_mask = 1'h1;
  assign ram_0_MPORT_40_en = reset;
  assign ram_0_MPORT_41_data = 1'h0;
  assign ram_0_MPORT_41_addr = 7'h29;
  assign ram_0_MPORT_41_mask = 1'h1;
  assign ram_0_MPORT_41_en = reset;
  assign ram_0_MPORT_42_data = 1'h0;
  assign ram_0_MPORT_42_addr = 7'h2a;
  assign ram_0_MPORT_42_mask = 1'h1;
  assign ram_0_MPORT_42_en = reset;
  assign ram_0_MPORT_43_data = 1'h0;
  assign ram_0_MPORT_43_addr = 7'h2b;
  assign ram_0_MPORT_43_mask = 1'h1;
  assign ram_0_MPORT_43_en = reset;
  assign ram_0_MPORT_44_data = 1'h0;
  assign ram_0_MPORT_44_addr = 7'h2c;
  assign ram_0_MPORT_44_mask = 1'h1;
  assign ram_0_MPORT_44_en = reset;
  assign ram_0_MPORT_45_data = 1'h0;
  assign ram_0_MPORT_45_addr = 7'h2d;
  assign ram_0_MPORT_45_mask = 1'h1;
  assign ram_0_MPORT_45_en = reset;
  assign ram_0_MPORT_46_data = 1'h0;
  assign ram_0_MPORT_46_addr = 7'h2e;
  assign ram_0_MPORT_46_mask = 1'h1;
  assign ram_0_MPORT_46_en = reset;
  assign ram_0_MPORT_47_data = 1'h0;
  assign ram_0_MPORT_47_addr = 7'h2f;
  assign ram_0_MPORT_47_mask = 1'h1;
  assign ram_0_MPORT_47_en = reset;
  assign ram_0_MPORT_48_data = 1'h0;
  assign ram_0_MPORT_48_addr = 7'h30;
  assign ram_0_MPORT_48_mask = 1'h1;
  assign ram_0_MPORT_48_en = reset;
  assign ram_0_MPORT_49_data = 1'h0;
  assign ram_0_MPORT_49_addr = 7'h31;
  assign ram_0_MPORT_49_mask = 1'h1;
  assign ram_0_MPORT_49_en = reset;
  assign ram_0_MPORT_50_data = 1'h0;
  assign ram_0_MPORT_50_addr = 7'h32;
  assign ram_0_MPORT_50_mask = 1'h1;
  assign ram_0_MPORT_50_en = reset;
  assign ram_0_MPORT_51_data = 1'h0;
  assign ram_0_MPORT_51_addr = 7'h33;
  assign ram_0_MPORT_51_mask = 1'h1;
  assign ram_0_MPORT_51_en = reset;
  assign ram_0_MPORT_52_data = 1'h0;
  assign ram_0_MPORT_52_addr = 7'h34;
  assign ram_0_MPORT_52_mask = 1'h1;
  assign ram_0_MPORT_52_en = reset;
  assign ram_0_MPORT_53_data = 1'h0;
  assign ram_0_MPORT_53_addr = 7'h35;
  assign ram_0_MPORT_53_mask = 1'h1;
  assign ram_0_MPORT_53_en = reset;
  assign ram_0_MPORT_54_data = 1'h0;
  assign ram_0_MPORT_54_addr = 7'h36;
  assign ram_0_MPORT_54_mask = 1'h1;
  assign ram_0_MPORT_54_en = reset;
  assign ram_0_MPORT_55_data = 1'h0;
  assign ram_0_MPORT_55_addr = 7'h37;
  assign ram_0_MPORT_55_mask = 1'h1;
  assign ram_0_MPORT_55_en = reset;
  assign ram_0_MPORT_56_data = 1'h0;
  assign ram_0_MPORT_56_addr = 7'h38;
  assign ram_0_MPORT_56_mask = 1'h1;
  assign ram_0_MPORT_56_en = reset;
  assign ram_0_MPORT_57_data = 1'h0;
  assign ram_0_MPORT_57_addr = 7'h39;
  assign ram_0_MPORT_57_mask = 1'h1;
  assign ram_0_MPORT_57_en = reset;
  assign ram_0_MPORT_58_data = 1'h0;
  assign ram_0_MPORT_58_addr = 7'h3a;
  assign ram_0_MPORT_58_mask = 1'h1;
  assign ram_0_MPORT_58_en = reset;
  assign ram_0_MPORT_59_data = 1'h0;
  assign ram_0_MPORT_59_addr = 7'h3b;
  assign ram_0_MPORT_59_mask = 1'h1;
  assign ram_0_MPORT_59_en = reset;
  assign ram_0_MPORT_60_data = 1'h0;
  assign ram_0_MPORT_60_addr = 7'h3c;
  assign ram_0_MPORT_60_mask = 1'h1;
  assign ram_0_MPORT_60_en = reset;
  assign ram_0_MPORT_61_data = 1'h0;
  assign ram_0_MPORT_61_addr = 7'h3d;
  assign ram_0_MPORT_61_mask = 1'h1;
  assign ram_0_MPORT_61_en = reset;
  assign ram_0_MPORT_62_data = 1'h0;
  assign ram_0_MPORT_62_addr = 7'h3e;
  assign ram_0_MPORT_62_mask = 1'h1;
  assign ram_0_MPORT_62_en = reset;
  assign ram_0_MPORT_63_data = 1'h0;
  assign ram_0_MPORT_63_addr = 7'h3f;
  assign ram_0_MPORT_63_mask = 1'h1;
  assign ram_0_MPORT_63_en = reset;
  assign ram_0_MPORT_64_data = 1'h0;
  assign ram_0_MPORT_64_addr = 7'h40;
  assign ram_0_MPORT_64_mask = 1'h1;
  assign ram_0_MPORT_64_en = reset;
  assign ram_0_MPORT_65_data = 1'h0;
  assign ram_0_MPORT_65_addr = 7'h41;
  assign ram_0_MPORT_65_mask = 1'h1;
  assign ram_0_MPORT_65_en = reset;
  assign ram_0_MPORT_66_data = 1'h0;
  assign ram_0_MPORT_66_addr = 7'h42;
  assign ram_0_MPORT_66_mask = 1'h1;
  assign ram_0_MPORT_66_en = reset;
  assign ram_0_MPORT_67_data = 1'h0;
  assign ram_0_MPORT_67_addr = 7'h43;
  assign ram_0_MPORT_67_mask = 1'h1;
  assign ram_0_MPORT_67_en = reset;
  assign ram_0_MPORT_68_data = 1'h0;
  assign ram_0_MPORT_68_addr = 7'h44;
  assign ram_0_MPORT_68_mask = 1'h1;
  assign ram_0_MPORT_68_en = reset;
  assign ram_0_MPORT_69_data = 1'h0;
  assign ram_0_MPORT_69_addr = 7'h45;
  assign ram_0_MPORT_69_mask = 1'h1;
  assign ram_0_MPORT_69_en = reset;
  assign ram_0_MPORT_70_data = 1'h0;
  assign ram_0_MPORT_70_addr = 7'h46;
  assign ram_0_MPORT_70_mask = 1'h1;
  assign ram_0_MPORT_70_en = reset;
  assign ram_0_MPORT_71_data = 1'h0;
  assign ram_0_MPORT_71_addr = 7'h47;
  assign ram_0_MPORT_71_mask = 1'h1;
  assign ram_0_MPORT_71_en = reset;
  assign ram_0_MPORT_72_data = 1'h0;
  assign ram_0_MPORT_72_addr = 7'h48;
  assign ram_0_MPORT_72_mask = 1'h1;
  assign ram_0_MPORT_72_en = reset;
  assign ram_0_MPORT_73_data = 1'h0;
  assign ram_0_MPORT_73_addr = 7'h49;
  assign ram_0_MPORT_73_mask = 1'h1;
  assign ram_0_MPORT_73_en = reset;
  assign ram_0_MPORT_74_data = 1'h0;
  assign ram_0_MPORT_74_addr = 7'h4a;
  assign ram_0_MPORT_74_mask = 1'h1;
  assign ram_0_MPORT_74_en = reset;
  assign ram_0_MPORT_75_data = 1'h0;
  assign ram_0_MPORT_75_addr = 7'h4b;
  assign ram_0_MPORT_75_mask = 1'h1;
  assign ram_0_MPORT_75_en = reset;
  assign ram_0_MPORT_76_data = 1'h0;
  assign ram_0_MPORT_76_addr = 7'h4c;
  assign ram_0_MPORT_76_mask = 1'h1;
  assign ram_0_MPORT_76_en = reset;
  assign ram_0_MPORT_77_data = 1'h0;
  assign ram_0_MPORT_77_addr = 7'h4d;
  assign ram_0_MPORT_77_mask = 1'h1;
  assign ram_0_MPORT_77_en = reset;
  assign ram_0_MPORT_78_data = 1'h0;
  assign ram_0_MPORT_78_addr = 7'h4e;
  assign ram_0_MPORT_78_mask = 1'h1;
  assign ram_0_MPORT_78_en = reset;
  assign ram_0_MPORT_79_data = 1'h0;
  assign ram_0_MPORT_79_addr = 7'h4f;
  assign ram_0_MPORT_79_mask = 1'h1;
  assign ram_0_MPORT_79_en = reset;
  assign ram_0_MPORT_80_data = 1'h0;
  assign ram_0_MPORT_80_addr = 7'h50;
  assign ram_0_MPORT_80_mask = 1'h1;
  assign ram_0_MPORT_80_en = reset;
  assign ram_0_MPORT_81_data = 1'h0;
  assign ram_0_MPORT_81_addr = 7'h51;
  assign ram_0_MPORT_81_mask = 1'h1;
  assign ram_0_MPORT_81_en = reset;
  assign ram_0_MPORT_82_data = 1'h0;
  assign ram_0_MPORT_82_addr = 7'h52;
  assign ram_0_MPORT_82_mask = 1'h1;
  assign ram_0_MPORT_82_en = reset;
  assign ram_0_MPORT_83_data = 1'h0;
  assign ram_0_MPORT_83_addr = 7'h53;
  assign ram_0_MPORT_83_mask = 1'h1;
  assign ram_0_MPORT_83_en = reset;
  assign ram_0_MPORT_84_data = 1'h0;
  assign ram_0_MPORT_84_addr = 7'h54;
  assign ram_0_MPORT_84_mask = 1'h1;
  assign ram_0_MPORT_84_en = reset;
  assign ram_0_MPORT_85_data = 1'h0;
  assign ram_0_MPORT_85_addr = 7'h55;
  assign ram_0_MPORT_85_mask = 1'h1;
  assign ram_0_MPORT_85_en = reset;
  assign ram_0_MPORT_86_data = 1'h0;
  assign ram_0_MPORT_86_addr = 7'h56;
  assign ram_0_MPORT_86_mask = 1'h1;
  assign ram_0_MPORT_86_en = reset;
  assign ram_0_MPORT_87_data = 1'h0;
  assign ram_0_MPORT_87_addr = 7'h57;
  assign ram_0_MPORT_87_mask = 1'h1;
  assign ram_0_MPORT_87_en = reset;
  assign ram_0_MPORT_88_data = 1'h0;
  assign ram_0_MPORT_88_addr = 7'h58;
  assign ram_0_MPORT_88_mask = 1'h1;
  assign ram_0_MPORT_88_en = reset;
  assign ram_0_MPORT_89_data = 1'h0;
  assign ram_0_MPORT_89_addr = 7'h59;
  assign ram_0_MPORT_89_mask = 1'h1;
  assign ram_0_MPORT_89_en = reset;
  assign ram_0_MPORT_90_data = 1'h0;
  assign ram_0_MPORT_90_addr = 7'h5a;
  assign ram_0_MPORT_90_mask = 1'h1;
  assign ram_0_MPORT_90_en = reset;
  assign ram_0_MPORT_91_data = 1'h0;
  assign ram_0_MPORT_91_addr = 7'h5b;
  assign ram_0_MPORT_91_mask = 1'h1;
  assign ram_0_MPORT_91_en = reset;
  assign ram_0_MPORT_92_data = 1'h0;
  assign ram_0_MPORT_92_addr = 7'h5c;
  assign ram_0_MPORT_92_mask = 1'h1;
  assign ram_0_MPORT_92_en = reset;
  assign ram_0_MPORT_93_data = 1'h0;
  assign ram_0_MPORT_93_addr = 7'h5d;
  assign ram_0_MPORT_93_mask = 1'h1;
  assign ram_0_MPORT_93_en = reset;
  assign ram_0_MPORT_94_data = 1'h0;
  assign ram_0_MPORT_94_addr = 7'h5e;
  assign ram_0_MPORT_94_mask = 1'h1;
  assign ram_0_MPORT_94_en = reset;
  assign ram_0_MPORT_95_data = 1'h0;
  assign ram_0_MPORT_95_addr = 7'h5f;
  assign ram_0_MPORT_95_mask = 1'h1;
  assign ram_0_MPORT_95_en = reset;
  assign ram_0_MPORT_96_data = 1'h0;
  assign ram_0_MPORT_96_addr = 7'h60;
  assign ram_0_MPORT_96_mask = 1'h1;
  assign ram_0_MPORT_96_en = reset;
  assign ram_0_MPORT_97_data = 1'h0;
  assign ram_0_MPORT_97_addr = 7'h61;
  assign ram_0_MPORT_97_mask = 1'h1;
  assign ram_0_MPORT_97_en = reset;
  assign ram_0_MPORT_98_data = 1'h0;
  assign ram_0_MPORT_98_addr = 7'h62;
  assign ram_0_MPORT_98_mask = 1'h1;
  assign ram_0_MPORT_98_en = reset;
  assign ram_0_MPORT_99_data = 1'h0;
  assign ram_0_MPORT_99_addr = 7'h63;
  assign ram_0_MPORT_99_mask = 1'h1;
  assign ram_0_MPORT_99_en = reset;
  assign ram_0_MPORT_100_data = 1'h0;
  assign ram_0_MPORT_100_addr = 7'h64;
  assign ram_0_MPORT_100_mask = 1'h1;
  assign ram_0_MPORT_100_en = reset;
  assign ram_0_MPORT_101_data = 1'h0;
  assign ram_0_MPORT_101_addr = 7'h65;
  assign ram_0_MPORT_101_mask = 1'h1;
  assign ram_0_MPORT_101_en = reset;
  assign ram_0_MPORT_102_data = 1'h0;
  assign ram_0_MPORT_102_addr = 7'h66;
  assign ram_0_MPORT_102_mask = 1'h1;
  assign ram_0_MPORT_102_en = reset;
  assign ram_0_MPORT_103_data = 1'h0;
  assign ram_0_MPORT_103_addr = 7'h67;
  assign ram_0_MPORT_103_mask = 1'h1;
  assign ram_0_MPORT_103_en = reset;
  assign ram_0_MPORT_104_data = 1'h0;
  assign ram_0_MPORT_104_addr = 7'h68;
  assign ram_0_MPORT_104_mask = 1'h1;
  assign ram_0_MPORT_104_en = reset;
  assign ram_0_MPORT_105_data = 1'h0;
  assign ram_0_MPORT_105_addr = 7'h69;
  assign ram_0_MPORT_105_mask = 1'h1;
  assign ram_0_MPORT_105_en = reset;
  assign ram_0_MPORT_106_data = 1'h0;
  assign ram_0_MPORT_106_addr = 7'h6a;
  assign ram_0_MPORT_106_mask = 1'h1;
  assign ram_0_MPORT_106_en = reset;
  assign ram_0_MPORT_107_data = 1'h0;
  assign ram_0_MPORT_107_addr = 7'h6b;
  assign ram_0_MPORT_107_mask = 1'h1;
  assign ram_0_MPORT_107_en = reset;
  assign ram_0_MPORT_108_data = 1'h0;
  assign ram_0_MPORT_108_addr = 7'h6c;
  assign ram_0_MPORT_108_mask = 1'h1;
  assign ram_0_MPORT_108_en = reset;
  assign ram_0_MPORT_109_data = 1'h0;
  assign ram_0_MPORT_109_addr = 7'h6d;
  assign ram_0_MPORT_109_mask = 1'h1;
  assign ram_0_MPORT_109_en = reset;
  assign ram_0_MPORT_110_data = 1'h0;
  assign ram_0_MPORT_110_addr = 7'h6e;
  assign ram_0_MPORT_110_mask = 1'h1;
  assign ram_0_MPORT_110_en = reset;
  assign ram_0_MPORT_111_data = 1'h0;
  assign ram_0_MPORT_111_addr = 7'h6f;
  assign ram_0_MPORT_111_mask = 1'h1;
  assign ram_0_MPORT_111_en = reset;
  assign ram_0_MPORT_112_data = 1'h0;
  assign ram_0_MPORT_112_addr = 7'h70;
  assign ram_0_MPORT_112_mask = 1'h1;
  assign ram_0_MPORT_112_en = reset;
  assign ram_0_MPORT_113_data = 1'h0;
  assign ram_0_MPORT_113_addr = 7'h71;
  assign ram_0_MPORT_113_mask = 1'h1;
  assign ram_0_MPORT_113_en = reset;
  assign ram_0_MPORT_114_data = 1'h0;
  assign ram_0_MPORT_114_addr = 7'h72;
  assign ram_0_MPORT_114_mask = 1'h1;
  assign ram_0_MPORT_114_en = reset;
  assign ram_0_MPORT_115_data = 1'h0;
  assign ram_0_MPORT_115_addr = 7'h73;
  assign ram_0_MPORT_115_mask = 1'h1;
  assign ram_0_MPORT_115_en = reset;
  assign ram_0_MPORT_116_data = 1'h0;
  assign ram_0_MPORT_116_addr = 7'h74;
  assign ram_0_MPORT_116_mask = 1'h1;
  assign ram_0_MPORT_116_en = reset;
  assign ram_0_MPORT_117_data = 1'h0;
  assign ram_0_MPORT_117_addr = 7'h75;
  assign ram_0_MPORT_117_mask = 1'h1;
  assign ram_0_MPORT_117_en = reset;
  assign ram_0_MPORT_118_data = 1'h0;
  assign ram_0_MPORT_118_addr = 7'h76;
  assign ram_0_MPORT_118_mask = 1'h1;
  assign ram_0_MPORT_118_en = reset;
  assign ram_0_MPORT_119_data = 1'h0;
  assign ram_0_MPORT_119_addr = 7'h77;
  assign ram_0_MPORT_119_mask = 1'h1;
  assign ram_0_MPORT_119_en = reset;
  assign ram_0_MPORT_120_data = 1'h0;
  assign ram_0_MPORT_120_addr = 7'h78;
  assign ram_0_MPORT_120_mask = 1'h1;
  assign ram_0_MPORT_120_en = reset;
  assign ram_0_MPORT_121_data = 1'h0;
  assign ram_0_MPORT_121_addr = 7'h79;
  assign ram_0_MPORT_121_mask = 1'h1;
  assign ram_0_MPORT_121_en = reset;
  assign ram_0_MPORT_122_data = 1'h0;
  assign ram_0_MPORT_122_addr = 7'h7a;
  assign ram_0_MPORT_122_mask = 1'h1;
  assign ram_0_MPORT_122_en = reset;
  assign ram_0_MPORT_123_data = 1'h0;
  assign ram_0_MPORT_123_addr = 7'h7b;
  assign ram_0_MPORT_123_mask = 1'h1;
  assign ram_0_MPORT_123_en = reset;
  assign ram_0_MPORT_124_data = 1'h0;
  assign ram_0_MPORT_124_addr = 7'h7c;
  assign ram_0_MPORT_124_mask = 1'h1;
  assign ram_0_MPORT_124_en = reset;
  assign ram_0_MPORT_125_data = 1'h0;
  assign ram_0_MPORT_125_addr = 7'h7d;
  assign ram_0_MPORT_125_mask = 1'h1;
  assign ram_0_MPORT_125_en = reset;
  assign ram_0_MPORT_126_data = 1'h0;
  assign ram_0_MPORT_126_addr = 7'h7e;
  assign ram_0_MPORT_126_mask = 1'h1;
  assign ram_0_MPORT_126_en = reset;
  assign ram_0_MPORT_127_data = 1'h0;
  assign ram_0_MPORT_127_addr = 7'h7f;
  assign ram_0_MPORT_127_mask = 1'h1;
  assign ram_0_MPORT_127_en = reset;
  assign ram_0_MPORT_128_data = 1'h1;
  assign ram_0_MPORT_128_addr = io_addr;
  assign ram_0_MPORT_128_mask = io_wmask[0];
  assign ram_0_MPORT_128_en = io_rw;
  assign ram_1_io_rdata_MPORT_en = ram_1_io_rdata_MPORT_en_pipe_0;
  assign ram_1_io_rdata_MPORT_addr = ram_1_io_rdata_MPORT_addr_pipe_0;
  assign ram_1_io_rdata_MPORT_data = ram_1[ram_1_io_rdata_MPORT_addr]; // @[SRAM.scala 36:26]
  assign ram_1_MPORT_data = 1'h0;
  assign ram_1_MPORT_addr = 7'h0;
  assign ram_1_MPORT_mask = 1'h1;
  assign ram_1_MPORT_en = reset;
  assign ram_1_MPORT_1_data = 1'h0;
  assign ram_1_MPORT_1_addr = 7'h1;
  assign ram_1_MPORT_1_mask = 1'h1;
  assign ram_1_MPORT_1_en = reset;
  assign ram_1_MPORT_2_data = 1'h0;
  assign ram_1_MPORT_2_addr = 7'h2;
  assign ram_1_MPORT_2_mask = 1'h1;
  assign ram_1_MPORT_2_en = reset;
  assign ram_1_MPORT_3_data = 1'h0;
  assign ram_1_MPORT_3_addr = 7'h3;
  assign ram_1_MPORT_3_mask = 1'h1;
  assign ram_1_MPORT_3_en = reset;
  assign ram_1_MPORT_4_data = 1'h0;
  assign ram_1_MPORT_4_addr = 7'h4;
  assign ram_1_MPORT_4_mask = 1'h1;
  assign ram_1_MPORT_4_en = reset;
  assign ram_1_MPORT_5_data = 1'h0;
  assign ram_1_MPORT_5_addr = 7'h5;
  assign ram_1_MPORT_5_mask = 1'h1;
  assign ram_1_MPORT_5_en = reset;
  assign ram_1_MPORT_6_data = 1'h0;
  assign ram_1_MPORT_6_addr = 7'h6;
  assign ram_1_MPORT_6_mask = 1'h1;
  assign ram_1_MPORT_6_en = reset;
  assign ram_1_MPORT_7_data = 1'h0;
  assign ram_1_MPORT_7_addr = 7'h7;
  assign ram_1_MPORT_7_mask = 1'h1;
  assign ram_1_MPORT_7_en = reset;
  assign ram_1_MPORT_8_data = 1'h0;
  assign ram_1_MPORT_8_addr = 7'h8;
  assign ram_1_MPORT_8_mask = 1'h1;
  assign ram_1_MPORT_8_en = reset;
  assign ram_1_MPORT_9_data = 1'h0;
  assign ram_1_MPORT_9_addr = 7'h9;
  assign ram_1_MPORT_9_mask = 1'h1;
  assign ram_1_MPORT_9_en = reset;
  assign ram_1_MPORT_10_data = 1'h0;
  assign ram_1_MPORT_10_addr = 7'ha;
  assign ram_1_MPORT_10_mask = 1'h1;
  assign ram_1_MPORT_10_en = reset;
  assign ram_1_MPORT_11_data = 1'h0;
  assign ram_1_MPORT_11_addr = 7'hb;
  assign ram_1_MPORT_11_mask = 1'h1;
  assign ram_1_MPORT_11_en = reset;
  assign ram_1_MPORT_12_data = 1'h0;
  assign ram_1_MPORT_12_addr = 7'hc;
  assign ram_1_MPORT_12_mask = 1'h1;
  assign ram_1_MPORT_12_en = reset;
  assign ram_1_MPORT_13_data = 1'h0;
  assign ram_1_MPORT_13_addr = 7'hd;
  assign ram_1_MPORT_13_mask = 1'h1;
  assign ram_1_MPORT_13_en = reset;
  assign ram_1_MPORT_14_data = 1'h0;
  assign ram_1_MPORT_14_addr = 7'he;
  assign ram_1_MPORT_14_mask = 1'h1;
  assign ram_1_MPORT_14_en = reset;
  assign ram_1_MPORT_15_data = 1'h0;
  assign ram_1_MPORT_15_addr = 7'hf;
  assign ram_1_MPORT_15_mask = 1'h1;
  assign ram_1_MPORT_15_en = reset;
  assign ram_1_MPORT_16_data = 1'h0;
  assign ram_1_MPORT_16_addr = 7'h10;
  assign ram_1_MPORT_16_mask = 1'h1;
  assign ram_1_MPORT_16_en = reset;
  assign ram_1_MPORT_17_data = 1'h0;
  assign ram_1_MPORT_17_addr = 7'h11;
  assign ram_1_MPORT_17_mask = 1'h1;
  assign ram_1_MPORT_17_en = reset;
  assign ram_1_MPORT_18_data = 1'h0;
  assign ram_1_MPORT_18_addr = 7'h12;
  assign ram_1_MPORT_18_mask = 1'h1;
  assign ram_1_MPORT_18_en = reset;
  assign ram_1_MPORT_19_data = 1'h0;
  assign ram_1_MPORT_19_addr = 7'h13;
  assign ram_1_MPORT_19_mask = 1'h1;
  assign ram_1_MPORT_19_en = reset;
  assign ram_1_MPORT_20_data = 1'h0;
  assign ram_1_MPORT_20_addr = 7'h14;
  assign ram_1_MPORT_20_mask = 1'h1;
  assign ram_1_MPORT_20_en = reset;
  assign ram_1_MPORT_21_data = 1'h0;
  assign ram_1_MPORT_21_addr = 7'h15;
  assign ram_1_MPORT_21_mask = 1'h1;
  assign ram_1_MPORT_21_en = reset;
  assign ram_1_MPORT_22_data = 1'h0;
  assign ram_1_MPORT_22_addr = 7'h16;
  assign ram_1_MPORT_22_mask = 1'h1;
  assign ram_1_MPORT_22_en = reset;
  assign ram_1_MPORT_23_data = 1'h0;
  assign ram_1_MPORT_23_addr = 7'h17;
  assign ram_1_MPORT_23_mask = 1'h1;
  assign ram_1_MPORT_23_en = reset;
  assign ram_1_MPORT_24_data = 1'h0;
  assign ram_1_MPORT_24_addr = 7'h18;
  assign ram_1_MPORT_24_mask = 1'h1;
  assign ram_1_MPORT_24_en = reset;
  assign ram_1_MPORT_25_data = 1'h0;
  assign ram_1_MPORT_25_addr = 7'h19;
  assign ram_1_MPORT_25_mask = 1'h1;
  assign ram_1_MPORT_25_en = reset;
  assign ram_1_MPORT_26_data = 1'h0;
  assign ram_1_MPORT_26_addr = 7'h1a;
  assign ram_1_MPORT_26_mask = 1'h1;
  assign ram_1_MPORT_26_en = reset;
  assign ram_1_MPORT_27_data = 1'h0;
  assign ram_1_MPORT_27_addr = 7'h1b;
  assign ram_1_MPORT_27_mask = 1'h1;
  assign ram_1_MPORT_27_en = reset;
  assign ram_1_MPORT_28_data = 1'h0;
  assign ram_1_MPORT_28_addr = 7'h1c;
  assign ram_1_MPORT_28_mask = 1'h1;
  assign ram_1_MPORT_28_en = reset;
  assign ram_1_MPORT_29_data = 1'h0;
  assign ram_1_MPORT_29_addr = 7'h1d;
  assign ram_1_MPORT_29_mask = 1'h1;
  assign ram_1_MPORT_29_en = reset;
  assign ram_1_MPORT_30_data = 1'h0;
  assign ram_1_MPORT_30_addr = 7'h1e;
  assign ram_1_MPORT_30_mask = 1'h1;
  assign ram_1_MPORT_30_en = reset;
  assign ram_1_MPORT_31_data = 1'h0;
  assign ram_1_MPORT_31_addr = 7'h1f;
  assign ram_1_MPORT_31_mask = 1'h1;
  assign ram_1_MPORT_31_en = reset;
  assign ram_1_MPORT_32_data = 1'h0;
  assign ram_1_MPORT_32_addr = 7'h20;
  assign ram_1_MPORT_32_mask = 1'h1;
  assign ram_1_MPORT_32_en = reset;
  assign ram_1_MPORT_33_data = 1'h0;
  assign ram_1_MPORT_33_addr = 7'h21;
  assign ram_1_MPORT_33_mask = 1'h1;
  assign ram_1_MPORT_33_en = reset;
  assign ram_1_MPORT_34_data = 1'h0;
  assign ram_1_MPORT_34_addr = 7'h22;
  assign ram_1_MPORT_34_mask = 1'h1;
  assign ram_1_MPORT_34_en = reset;
  assign ram_1_MPORT_35_data = 1'h0;
  assign ram_1_MPORT_35_addr = 7'h23;
  assign ram_1_MPORT_35_mask = 1'h1;
  assign ram_1_MPORT_35_en = reset;
  assign ram_1_MPORT_36_data = 1'h0;
  assign ram_1_MPORT_36_addr = 7'h24;
  assign ram_1_MPORT_36_mask = 1'h1;
  assign ram_1_MPORT_36_en = reset;
  assign ram_1_MPORT_37_data = 1'h0;
  assign ram_1_MPORT_37_addr = 7'h25;
  assign ram_1_MPORT_37_mask = 1'h1;
  assign ram_1_MPORT_37_en = reset;
  assign ram_1_MPORT_38_data = 1'h0;
  assign ram_1_MPORT_38_addr = 7'h26;
  assign ram_1_MPORT_38_mask = 1'h1;
  assign ram_1_MPORT_38_en = reset;
  assign ram_1_MPORT_39_data = 1'h0;
  assign ram_1_MPORT_39_addr = 7'h27;
  assign ram_1_MPORT_39_mask = 1'h1;
  assign ram_1_MPORT_39_en = reset;
  assign ram_1_MPORT_40_data = 1'h0;
  assign ram_1_MPORT_40_addr = 7'h28;
  assign ram_1_MPORT_40_mask = 1'h1;
  assign ram_1_MPORT_40_en = reset;
  assign ram_1_MPORT_41_data = 1'h0;
  assign ram_1_MPORT_41_addr = 7'h29;
  assign ram_1_MPORT_41_mask = 1'h1;
  assign ram_1_MPORT_41_en = reset;
  assign ram_1_MPORT_42_data = 1'h0;
  assign ram_1_MPORT_42_addr = 7'h2a;
  assign ram_1_MPORT_42_mask = 1'h1;
  assign ram_1_MPORT_42_en = reset;
  assign ram_1_MPORT_43_data = 1'h0;
  assign ram_1_MPORT_43_addr = 7'h2b;
  assign ram_1_MPORT_43_mask = 1'h1;
  assign ram_1_MPORT_43_en = reset;
  assign ram_1_MPORT_44_data = 1'h0;
  assign ram_1_MPORT_44_addr = 7'h2c;
  assign ram_1_MPORT_44_mask = 1'h1;
  assign ram_1_MPORT_44_en = reset;
  assign ram_1_MPORT_45_data = 1'h0;
  assign ram_1_MPORT_45_addr = 7'h2d;
  assign ram_1_MPORT_45_mask = 1'h1;
  assign ram_1_MPORT_45_en = reset;
  assign ram_1_MPORT_46_data = 1'h0;
  assign ram_1_MPORT_46_addr = 7'h2e;
  assign ram_1_MPORT_46_mask = 1'h1;
  assign ram_1_MPORT_46_en = reset;
  assign ram_1_MPORT_47_data = 1'h0;
  assign ram_1_MPORT_47_addr = 7'h2f;
  assign ram_1_MPORT_47_mask = 1'h1;
  assign ram_1_MPORT_47_en = reset;
  assign ram_1_MPORT_48_data = 1'h0;
  assign ram_1_MPORT_48_addr = 7'h30;
  assign ram_1_MPORT_48_mask = 1'h1;
  assign ram_1_MPORT_48_en = reset;
  assign ram_1_MPORT_49_data = 1'h0;
  assign ram_1_MPORT_49_addr = 7'h31;
  assign ram_1_MPORT_49_mask = 1'h1;
  assign ram_1_MPORT_49_en = reset;
  assign ram_1_MPORT_50_data = 1'h0;
  assign ram_1_MPORT_50_addr = 7'h32;
  assign ram_1_MPORT_50_mask = 1'h1;
  assign ram_1_MPORT_50_en = reset;
  assign ram_1_MPORT_51_data = 1'h0;
  assign ram_1_MPORT_51_addr = 7'h33;
  assign ram_1_MPORT_51_mask = 1'h1;
  assign ram_1_MPORT_51_en = reset;
  assign ram_1_MPORT_52_data = 1'h0;
  assign ram_1_MPORT_52_addr = 7'h34;
  assign ram_1_MPORT_52_mask = 1'h1;
  assign ram_1_MPORT_52_en = reset;
  assign ram_1_MPORT_53_data = 1'h0;
  assign ram_1_MPORT_53_addr = 7'h35;
  assign ram_1_MPORT_53_mask = 1'h1;
  assign ram_1_MPORT_53_en = reset;
  assign ram_1_MPORT_54_data = 1'h0;
  assign ram_1_MPORT_54_addr = 7'h36;
  assign ram_1_MPORT_54_mask = 1'h1;
  assign ram_1_MPORT_54_en = reset;
  assign ram_1_MPORT_55_data = 1'h0;
  assign ram_1_MPORT_55_addr = 7'h37;
  assign ram_1_MPORT_55_mask = 1'h1;
  assign ram_1_MPORT_55_en = reset;
  assign ram_1_MPORT_56_data = 1'h0;
  assign ram_1_MPORT_56_addr = 7'h38;
  assign ram_1_MPORT_56_mask = 1'h1;
  assign ram_1_MPORT_56_en = reset;
  assign ram_1_MPORT_57_data = 1'h0;
  assign ram_1_MPORT_57_addr = 7'h39;
  assign ram_1_MPORT_57_mask = 1'h1;
  assign ram_1_MPORT_57_en = reset;
  assign ram_1_MPORT_58_data = 1'h0;
  assign ram_1_MPORT_58_addr = 7'h3a;
  assign ram_1_MPORT_58_mask = 1'h1;
  assign ram_1_MPORT_58_en = reset;
  assign ram_1_MPORT_59_data = 1'h0;
  assign ram_1_MPORT_59_addr = 7'h3b;
  assign ram_1_MPORT_59_mask = 1'h1;
  assign ram_1_MPORT_59_en = reset;
  assign ram_1_MPORT_60_data = 1'h0;
  assign ram_1_MPORT_60_addr = 7'h3c;
  assign ram_1_MPORT_60_mask = 1'h1;
  assign ram_1_MPORT_60_en = reset;
  assign ram_1_MPORT_61_data = 1'h0;
  assign ram_1_MPORT_61_addr = 7'h3d;
  assign ram_1_MPORT_61_mask = 1'h1;
  assign ram_1_MPORT_61_en = reset;
  assign ram_1_MPORT_62_data = 1'h0;
  assign ram_1_MPORT_62_addr = 7'h3e;
  assign ram_1_MPORT_62_mask = 1'h1;
  assign ram_1_MPORT_62_en = reset;
  assign ram_1_MPORT_63_data = 1'h0;
  assign ram_1_MPORT_63_addr = 7'h3f;
  assign ram_1_MPORT_63_mask = 1'h1;
  assign ram_1_MPORT_63_en = reset;
  assign ram_1_MPORT_64_data = 1'h0;
  assign ram_1_MPORT_64_addr = 7'h40;
  assign ram_1_MPORT_64_mask = 1'h1;
  assign ram_1_MPORT_64_en = reset;
  assign ram_1_MPORT_65_data = 1'h0;
  assign ram_1_MPORT_65_addr = 7'h41;
  assign ram_1_MPORT_65_mask = 1'h1;
  assign ram_1_MPORT_65_en = reset;
  assign ram_1_MPORT_66_data = 1'h0;
  assign ram_1_MPORT_66_addr = 7'h42;
  assign ram_1_MPORT_66_mask = 1'h1;
  assign ram_1_MPORT_66_en = reset;
  assign ram_1_MPORT_67_data = 1'h0;
  assign ram_1_MPORT_67_addr = 7'h43;
  assign ram_1_MPORT_67_mask = 1'h1;
  assign ram_1_MPORT_67_en = reset;
  assign ram_1_MPORT_68_data = 1'h0;
  assign ram_1_MPORT_68_addr = 7'h44;
  assign ram_1_MPORT_68_mask = 1'h1;
  assign ram_1_MPORT_68_en = reset;
  assign ram_1_MPORT_69_data = 1'h0;
  assign ram_1_MPORT_69_addr = 7'h45;
  assign ram_1_MPORT_69_mask = 1'h1;
  assign ram_1_MPORT_69_en = reset;
  assign ram_1_MPORT_70_data = 1'h0;
  assign ram_1_MPORT_70_addr = 7'h46;
  assign ram_1_MPORT_70_mask = 1'h1;
  assign ram_1_MPORT_70_en = reset;
  assign ram_1_MPORT_71_data = 1'h0;
  assign ram_1_MPORT_71_addr = 7'h47;
  assign ram_1_MPORT_71_mask = 1'h1;
  assign ram_1_MPORT_71_en = reset;
  assign ram_1_MPORT_72_data = 1'h0;
  assign ram_1_MPORT_72_addr = 7'h48;
  assign ram_1_MPORT_72_mask = 1'h1;
  assign ram_1_MPORT_72_en = reset;
  assign ram_1_MPORT_73_data = 1'h0;
  assign ram_1_MPORT_73_addr = 7'h49;
  assign ram_1_MPORT_73_mask = 1'h1;
  assign ram_1_MPORT_73_en = reset;
  assign ram_1_MPORT_74_data = 1'h0;
  assign ram_1_MPORT_74_addr = 7'h4a;
  assign ram_1_MPORT_74_mask = 1'h1;
  assign ram_1_MPORT_74_en = reset;
  assign ram_1_MPORT_75_data = 1'h0;
  assign ram_1_MPORT_75_addr = 7'h4b;
  assign ram_1_MPORT_75_mask = 1'h1;
  assign ram_1_MPORT_75_en = reset;
  assign ram_1_MPORT_76_data = 1'h0;
  assign ram_1_MPORT_76_addr = 7'h4c;
  assign ram_1_MPORT_76_mask = 1'h1;
  assign ram_1_MPORT_76_en = reset;
  assign ram_1_MPORT_77_data = 1'h0;
  assign ram_1_MPORT_77_addr = 7'h4d;
  assign ram_1_MPORT_77_mask = 1'h1;
  assign ram_1_MPORT_77_en = reset;
  assign ram_1_MPORT_78_data = 1'h0;
  assign ram_1_MPORT_78_addr = 7'h4e;
  assign ram_1_MPORT_78_mask = 1'h1;
  assign ram_1_MPORT_78_en = reset;
  assign ram_1_MPORT_79_data = 1'h0;
  assign ram_1_MPORT_79_addr = 7'h4f;
  assign ram_1_MPORT_79_mask = 1'h1;
  assign ram_1_MPORT_79_en = reset;
  assign ram_1_MPORT_80_data = 1'h0;
  assign ram_1_MPORT_80_addr = 7'h50;
  assign ram_1_MPORT_80_mask = 1'h1;
  assign ram_1_MPORT_80_en = reset;
  assign ram_1_MPORT_81_data = 1'h0;
  assign ram_1_MPORT_81_addr = 7'h51;
  assign ram_1_MPORT_81_mask = 1'h1;
  assign ram_1_MPORT_81_en = reset;
  assign ram_1_MPORT_82_data = 1'h0;
  assign ram_1_MPORT_82_addr = 7'h52;
  assign ram_1_MPORT_82_mask = 1'h1;
  assign ram_1_MPORT_82_en = reset;
  assign ram_1_MPORT_83_data = 1'h0;
  assign ram_1_MPORT_83_addr = 7'h53;
  assign ram_1_MPORT_83_mask = 1'h1;
  assign ram_1_MPORT_83_en = reset;
  assign ram_1_MPORT_84_data = 1'h0;
  assign ram_1_MPORT_84_addr = 7'h54;
  assign ram_1_MPORT_84_mask = 1'h1;
  assign ram_1_MPORT_84_en = reset;
  assign ram_1_MPORT_85_data = 1'h0;
  assign ram_1_MPORT_85_addr = 7'h55;
  assign ram_1_MPORT_85_mask = 1'h1;
  assign ram_1_MPORT_85_en = reset;
  assign ram_1_MPORT_86_data = 1'h0;
  assign ram_1_MPORT_86_addr = 7'h56;
  assign ram_1_MPORT_86_mask = 1'h1;
  assign ram_1_MPORT_86_en = reset;
  assign ram_1_MPORT_87_data = 1'h0;
  assign ram_1_MPORT_87_addr = 7'h57;
  assign ram_1_MPORT_87_mask = 1'h1;
  assign ram_1_MPORT_87_en = reset;
  assign ram_1_MPORT_88_data = 1'h0;
  assign ram_1_MPORT_88_addr = 7'h58;
  assign ram_1_MPORT_88_mask = 1'h1;
  assign ram_1_MPORT_88_en = reset;
  assign ram_1_MPORT_89_data = 1'h0;
  assign ram_1_MPORT_89_addr = 7'h59;
  assign ram_1_MPORT_89_mask = 1'h1;
  assign ram_1_MPORT_89_en = reset;
  assign ram_1_MPORT_90_data = 1'h0;
  assign ram_1_MPORT_90_addr = 7'h5a;
  assign ram_1_MPORT_90_mask = 1'h1;
  assign ram_1_MPORT_90_en = reset;
  assign ram_1_MPORT_91_data = 1'h0;
  assign ram_1_MPORT_91_addr = 7'h5b;
  assign ram_1_MPORT_91_mask = 1'h1;
  assign ram_1_MPORT_91_en = reset;
  assign ram_1_MPORT_92_data = 1'h0;
  assign ram_1_MPORT_92_addr = 7'h5c;
  assign ram_1_MPORT_92_mask = 1'h1;
  assign ram_1_MPORT_92_en = reset;
  assign ram_1_MPORT_93_data = 1'h0;
  assign ram_1_MPORT_93_addr = 7'h5d;
  assign ram_1_MPORT_93_mask = 1'h1;
  assign ram_1_MPORT_93_en = reset;
  assign ram_1_MPORT_94_data = 1'h0;
  assign ram_1_MPORT_94_addr = 7'h5e;
  assign ram_1_MPORT_94_mask = 1'h1;
  assign ram_1_MPORT_94_en = reset;
  assign ram_1_MPORT_95_data = 1'h0;
  assign ram_1_MPORT_95_addr = 7'h5f;
  assign ram_1_MPORT_95_mask = 1'h1;
  assign ram_1_MPORT_95_en = reset;
  assign ram_1_MPORT_96_data = 1'h0;
  assign ram_1_MPORT_96_addr = 7'h60;
  assign ram_1_MPORT_96_mask = 1'h1;
  assign ram_1_MPORT_96_en = reset;
  assign ram_1_MPORT_97_data = 1'h0;
  assign ram_1_MPORT_97_addr = 7'h61;
  assign ram_1_MPORT_97_mask = 1'h1;
  assign ram_1_MPORT_97_en = reset;
  assign ram_1_MPORT_98_data = 1'h0;
  assign ram_1_MPORT_98_addr = 7'h62;
  assign ram_1_MPORT_98_mask = 1'h1;
  assign ram_1_MPORT_98_en = reset;
  assign ram_1_MPORT_99_data = 1'h0;
  assign ram_1_MPORT_99_addr = 7'h63;
  assign ram_1_MPORT_99_mask = 1'h1;
  assign ram_1_MPORT_99_en = reset;
  assign ram_1_MPORT_100_data = 1'h0;
  assign ram_1_MPORT_100_addr = 7'h64;
  assign ram_1_MPORT_100_mask = 1'h1;
  assign ram_1_MPORT_100_en = reset;
  assign ram_1_MPORT_101_data = 1'h0;
  assign ram_1_MPORT_101_addr = 7'h65;
  assign ram_1_MPORT_101_mask = 1'h1;
  assign ram_1_MPORT_101_en = reset;
  assign ram_1_MPORT_102_data = 1'h0;
  assign ram_1_MPORT_102_addr = 7'h66;
  assign ram_1_MPORT_102_mask = 1'h1;
  assign ram_1_MPORT_102_en = reset;
  assign ram_1_MPORT_103_data = 1'h0;
  assign ram_1_MPORT_103_addr = 7'h67;
  assign ram_1_MPORT_103_mask = 1'h1;
  assign ram_1_MPORT_103_en = reset;
  assign ram_1_MPORT_104_data = 1'h0;
  assign ram_1_MPORT_104_addr = 7'h68;
  assign ram_1_MPORT_104_mask = 1'h1;
  assign ram_1_MPORT_104_en = reset;
  assign ram_1_MPORT_105_data = 1'h0;
  assign ram_1_MPORT_105_addr = 7'h69;
  assign ram_1_MPORT_105_mask = 1'h1;
  assign ram_1_MPORT_105_en = reset;
  assign ram_1_MPORT_106_data = 1'h0;
  assign ram_1_MPORT_106_addr = 7'h6a;
  assign ram_1_MPORT_106_mask = 1'h1;
  assign ram_1_MPORT_106_en = reset;
  assign ram_1_MPORT_107_data = 1'h0;
  assign ram_1_MPORT_107_addr = 7'h6b;
  assign ram_1_MPORT_107_mask = 1'h1;
  assign ram_1_MPORT_107_en = reset;
  assign ram_1_MPORT_108_data = 1'h0;
  assign ram_1_MPORT_108_addr = 7'h6c;
  assign ram_1_MPORT_108_mask = 1'h1;
  assign ram_1_MPORT_108_en = reset;
  assign ram_1_MPORT_109_data = 1'h0;
  assign ram_1_MPORT_109_addr = 7'h6d;
  assign ram_1_MPORT_109_mask = 1'h1;
  assign ram_1_MPORT_109_en = reset;
  assign ram_1_MPORT_110_data = 1'h0;
  assign ram_1_MPORT_110_addr = 7'h6e;
  assign ram_1_MPORT_110_mask = 1'h1;
  assign ram_1_MPORT_110_en = reset;
  assign ram_1_MPORT_111_data = 1'h0;
  assign ram_1_MPORT_111_addr = 7'h6f;
  assign ram_1_MPORT_111_mask = 1'h1;
  assign ram_1_MPORT_111_en = reset;
  assign ram_1_MPORT_112_data = 1'h0;
  assign ram_1_MPORT_112_addr = 7'h70;
  assign ram_1_MPORT_112_mask = 1'h1;
  assign ram_1_MPORT_112_en = reset;
  assign ram_1_MPORT_113_data = 1'h0;
  assign ram_1_MPORT_113_addr = 7'h71;
  assign ram_1_MPORT_113_mask = 1'h1;
  assign ram_1_MPORT_113_en = reset;
  assign ram_1_MPORT_114_data = 1'h0;
  assign ram_1_MPORT_114_addr = 7'h72;
  assign ram_1_MPORT_114_mask = 1'h1;
  assign ram_1_MPORT_114_en = reset;
  assign ram_1_MPORT_115_data = 1'h0;
  assign ram_1_MPORT_115_addr = 7'h73;
  assign ram_1_MPORT_115_mask = 1'h1;
  assign ram_1_MPORT_115_en = reset;
  assign ram_1_MPORT_116_data = 1'h0;
  assign ram_1_MPORT_116_addr = 7'h74;
  assign ram_1_MPORT_116_mask = 1'h1;
  assign ram_1_MPORT_116_en = reset;
  assign ram_1_MPORT_117_data = 1'h0;
  assign ram_1_MPORT_117_addr = 7'h75;
  assign ram_1_MPORT_117_mask = 1'h1;
  assign ram_1_MPORT_117_en = reset;
  assign ram_1_MPORT_118_data = 1'h0;
  assign ram_1_MPORT_118_addr = 7'h76;
  assign ram_1_MPORT_118_mask = 1'h1;
  assign ram_1_MPORT_118_en = reset;
  assign ram_1_MPORT_119_data = 1'h0;
  assign ram_1_MPORT_119_addr = 7'h77;
  assign ram_1_MPORT_119_mask = 1'h1;
  assign ram_1_MPORT_119_en = reset;
  assign ram_1_MPORT_120_data = 1'h0;
  assign ram_1_MPORT_120_addr = 7'h78;
  assign ram_1_MPORT_120_mask = 1'h1;
  assign ram_1_MPORT_120_en = reset;
  assign ram_1_MPORT_121_data = 1'h0;
  assign ram_1_MPORT_121_addr = 7'h79;
  assign ram_1_MPORT_121_mask = 1'h1;
  assign ram_1_MPORT_121_en = reset;
  assign ram_1_MPORT_122_data = 1'h0;
  assign ram_1_MPORT_122_addr = 7'h7a;
  assign ram_1_MPORT_122_mask = 1'h1;
  assign ram_1_MPORT_122_en = reset;
  assign ram_1_MPORT_123_data = 1'h0;
  assign ram_1_MPORT_123_addr = 7'h7b;
  assign ram_1_MPORT_123_mask = 1'h1;
  assign ram_1_MPORT_123_en = reset;
  assign ram_1_MPORT_124_data = 1'h0;
  assign ram_1_MPORT_124_addr = 7'h7c;
  assign ram_1_MPORT_124_mask = 1'h1;
  assign ram_1_MPORT_124_en = reset;
  assign ram_1_MPORT_125_data = 1'h0;
  assign ram_1_MPORT_125_addr = 7'h7d;
  assign ram_1_MPORT_125_mask = 1'h1;
  assign ram_1_MPORT_125_en = reset;
  assign ram_1_MPORT_126_data = 1'h0;
  assign ram_1_MPORT_126_addr = 7'h7e;
  assign ram_1_MPORT_126_mask = 1'h1;
  assign ram_1_MPORT_126_en = reset;
  assign ram_1_MPORT_127_data = 1'h0;
  assign ram_1_MPORT_127_addr = 7'h7f;
  assign ram_1_MPORT_127_mask = 1'h1;
  assign ram_1_MPORT_127_en = reset;
  assign ram_1_MPORT_128_data = 1'h1;
  assign ram_1_MPORT_128_addr = io_addr;
  assign ram_1_MPORT_128_mask = io_wmask[1];
  assign ram_1_MPORT_128_en = io_rw;
  assign ram_2_io_rdata_MPORT_en = ram_2_io_rdata_MPORT_en_pipe_0;
  assign ram_2_io_rdata_MPORT_addr = ram_2_io_rdata_MPORT_addr_pipe_0;
  assign ram_2_io_rdata_MPORT_data = ram_2[ram_2_io_rdata_MPORT_addr]; // @[SRAM.scala 36:26]
  assign ram_2_MPORT_data = 1'h0;
  assign ram_2_MPORT_addr = 7'h0;
  assign ram_2_MPORT_mask = 1'h1;
  assign ram_2_MPORT_en = reset;
  assign ram_2_MPORT_1_data = 1'h0;
  assign ram_2_MPORT_1_addr = 7'h1;
  assign ram_2_MPORT_1_mask = 1'h1;
  assign ram_2_MPORT_1_en = reset;
  assign ram_2_MPORT_2_data = 1'h0;
  assign ram_2_MPORT_2_addr = 7'h2;
  assign ram_2_MPORT_2_mask = 1'h1;
  assign ram_2_MPORT_2_en = reset;
  assign ram_2_MPORT_3_data = 1'h0;
  assign ram_2_MPORT_3_addr = 7'h3;
  assign ram_2_MPORT_3_mask = 1'h1;
  assign ram_2_MPORT_3_en = reset;
  assign ram_2_MPORT_4_data = 1'h0;
  assign ram_2_MPORT_4_addr = 7'h4;
  assign ram_2_MPORT_4_mask = 1'h1;
  assign ram_2_MPORT_4_en = reset;
  assign ram_2_MPORT_5_data = 1'h0;
  assign ram_2_MPORT_5_addr = 7'h5;
  assign ram_2_MPORT_5_mask = 1'h1;
  assign ram_2_MPORT_5_en = reset;
  assign ram_2_MPORT_6_data = 1'h0;
  assign ram_2_MPORT_6_addr = 7'h6;
  assign ram_2_MPORT_6_mask = 1'h1;
  assign ram_2_MPORT_6_en = reset;
  assign ram_2_MPORT_7_data = 1'h0;
  assign ram_2_MPORT_7_addr = 7'h7;
  assign ram_2_MPORT_7_mask = 1'h1;
  assign ram_2_MPORT_7_en = reset;
  assign ram_2_MPORT_8_data = 1'h0;
  assign ram_2_MPORT_8_addr = 7'h8;
  assign ram_2_MPORT_8_mask = 1'h1;
  assign ram_2_MPORT_8_en = reset;
  assign ram_2_MPORT_9_data = 1'h0;
  assign ram_2_MPORT_9_addr = 7'h9;
  assign ram_2_MPORT_9_mask = 1'h1;
  assign ram_2_MPORT_9_en = reset;
  assign ram_2_MPORT_10_data = 1'h0;
  assign ram_2_MPORT_10_addr = 7'ha;
  assign ram_2_MPORT_10_mask = 1'h1;
  assign ram_2_MPORT_10_en = reset;
  assign ram_2_MPORT_11_data = 1'h0;
  assign ram_2_MPORT_11_addr = 7'hb;
  assign ram_2_MPORT_11_mask = 1'h1;
  assign ram_2_MPORT_11_en = reset;
  assign ram_2_MPORT_12_data = 1'h0;
  assign ram_2_MPORT_12_addr = 7'hc;
  assign ram_2_MPORT_12_mask = 1'h1;
  assign ram_2_MPORT_12_en = reset;
  assign ram_2_MPORT_13_data = 1'h0;
  assign ram_2_MPORT_13_addr = 7'hd;
  assign ram_2_MPORT_13_mask = 1'h1;
  assign ram_2_MPORT_13_en = reset;
  assign ram_2_MPORT_14_data = 1'h0;
  assign ram_2_MPORT_14_addr = 7'he;
  assign ram_2_MPORT_14_mask = 1'h1;
  assign ram_2_MPORT_14_en = reset;
  assign ram_2_MPORT_15_data = 1'h0;
  assign ram_2_MPORT_15_addr = 7'hf;
  assign ram_2_MPORT_15_mask = 1'h1;
  assign ram_2_MPORT_15_en = reset;
  assign ram_2_MPORT_16_data = 1'h0;
  assign ram_2_MPORT_16_addr = 7'h10;
  assign ram_2_MPORT_16_mask = 1'h1;
  assign ram_2_MPORT_16_en = reset;
  assign ram_2_MPORT_17_data = 1'h0;
  assign ram_2_MPORT_17_addr = 7'h11;
  assign ram_2_MPORT_17_mask = 1'h1;
  assign ram_2_MPORT_17_en = reset;
  assign ram_2_MPORT_18_data = 1'h0;
  assign ram_2_MPORT_18_addr = 7'h12;
  assign ram_2_MPORT_18_mask = 1'h1;
  assign ram_2_MPORT_18_en = reset;
  assign ram_2_MPORT_19_data = 1'h0;
  assign ram_2_MPORT_19_addr = 7'h13;
  assign ram_2_MPORT_19_mask = 1'h1;
  assign ram_2_MPORT_19_en = reset;
  assign ram_2_MPORT_20_data = 1'h0;
  assign ram_2_MPORT_20_addr = 7'h14;
  assign ram_2_MPORT_20_mask = 1'h1;
  assign ram_2_MPORT_20_en = reset;
  assign ram_2_MPORT_21_data = 1'h0;
  assign ram_2_MPORT_21_addr = 7'h15;
  assign ram_2_MPORT_21_mask = 1'h1;
  assign ram_2_MPORT_21_en = reset;
  assign ram_2_MPORT_22_data = 1'h0;
  assign ram_2_MPORT_22_addr = 7'h16;
  assign ram_2_MPORT_22_mask = 1'h1;
  assign ram_2_MPORT_22_en = reset;
  assign ram_2_MPORT_23_data = 1'h0;
  assign ram_2_MPORT_23_addr = 7'h17;
  assign ram_2_MPORT_23_mask = 1'h1;
  assign ram_2_MPORT_23_en = reset;
  assign ram_2_MPORT_24_data = 1'h0;
  assign ram_2_MPORT_24_addr = 7'h18;
  assign ram_2_MPORT_24_mask = 1'h1;
  assign ram_2_MPORT_24_en = reset;
  assign ram_2_MPORT_25_data = 1'h0;
  assign ram_2_MPORT_25_addr = 7'h19;
  assign ram_2_MPORT_25_mask = 1'h1;
  assign ram_2_MPORT_25_en = reset;
  assign ram_2_MPORT_26_data = 1'h0;
  assign ram_2_MPORT_26_addr = 7'h1a;
  assign ram_2_MPORT_26_mask = 1'h1;
  assign ram_2_MPORT_26_en = reset;
  assign ram_2_MPORT_27_data = 1'h0;
  assign ram_2_MPORT_27_addr = 7'h1b;
  assign ram_2_MPORT_27_mask = 1'h1;
  assign ram_2_MPORT_27_en = reset;
  assign ram_2_MPORT_28_data = 1'h0;
  assign ram_2_MPORT_28_addr = 7'h1c;
  assign ram_2_MPORT_28_mask = 1'h1;
  assign ram_2_MPORT_28_en = reset;
  assign ram_2_MPORT_29_data = 1'h0;
  assign ram_2_MPORT_29_addr = 7'h1d;
  assign ram_2_MPORT_29_mask = 1'h1;
  assign ram_2_MPORT_29_en = reset;
  assign ram_2_MPORT_30_data = 1'h0;
  assign ram_2_MPORT_30_addr = 7'h1e;
  assign ram_2_MPORT_30_mask = 1'h1;
  assign ram_2_MPORT_30_en = reset;
  assign ram_2_MPORT_31_data = 1'h0;
  assign ram_2_MPORT_31_addr = 7'h1f;
  assign ram_2_MPORT_31_mask = 1'h1;
  assign ram_2_MPORT_31_en = reset;
  assign ram_2_MPORT_32_data = 1'h0;
  assign ram_2_MPORT_32_addr = 7'h20;
  assign ram_2_MPORT_32_mask = 1'h1;
  assign ram_2_MPORT_32_en = reset;
  assign ram_2_MPORT_33_data = 1'h0;
  assign ram_2_MPORT_33_addr = 7'h21;
  assign ram_2_MPORT_33_mask = 1'h1;
  assign ram_2_MPORT_33_en = reset;
  assign ram_2_MPORT_34_data = 1'h0;
  assign ram_2_MPORT_34_addr = 7'h22;
  assign ram_2_MPORT_34_mask = 1'h1;
  assign ram_2_MPORT_34_en = reset;
  assign ram_2_MPORT_35_data = 1'h0;
  assign ram_2_MPORT_35_addr = 7'h23;
  assign ram_2_MPORT_35_mask = 1'h1;
  assign ram_2_MPORT_35_en = reset;
  assign ram_2_MPORT_36_data = 1'h0;
  assign ram_2_MPORT_36_addr = 7'h24;
  assign ram_2_MPORT_36_mask = 1'h1;
  assign ram_2_MPORT_36_en = reset;
  assign ram_2_MPORT_37_data = 1'h0;
  assign ram_2_MPORT_37_addr = 7'h25;
  assign ram_2_MPORT_37_mask = 1'h1;
  assign ram_2_MPORT_37_en = reset;
  assign ram_2_MPORT_38_data = 1'h0;
  assign ram_2_MPORT_38_addr = 7'h26;
  assign ram_2_MPORT_38_mask = 1'h1;
  assign ram_2_MPORT_38_en = reset;
  assign ram_2_MPORT_39_data = 1'h0;
  assign ram_2_MPORT_39_addr = 7'h27;
  assign ram_2_MPORT_39_mask = 1'h1;
  assign ram_2_MPORT_39_en = reset;
  assign ram_2_MPORT_40_data = 1'h0;
  assign ram_2_MPORT_40_addr = 7'h28;
  assign ram_2_MPORT_40_mask = 1'h1;
  assign ram_2_MPORT_40_en = reset;
  assign ram_2_MPORT_41_data = 1'h0;
  assign ram_2_MPORT_41_addr = 7'h29;
  assign ram_2_MPORT_41_mask = 1'h1;
  assign ram_2_MPORT_41_en = reset;
  assign ram_2_MPORT_42_data = 1'h0;
  assign ram_2_MPORT_42_addr = 7'h2a;
  assign ram_2_MPORT_42_mask = 1'h1;
  assign ram_2_MPORT_42_en = reset;
  assign ram_2_MPORT_43_data = 1'h0;
  assign ram_2_MPORT_43_addr = 7'h2b;
  assign ram_2_MPORT_43_mask = 1'h1;
  assign ram_2_MPORT_43_en = reset;
  assign ram_2_MPORT_44_data = 1'h0;
  assign ram_2_MPORT_44_addr = 7'h2c;
  assign ram_2_MPORT_44_mask = 1'h1;
  assign ram_2_MPORT_44_en = reset;
  assign ram_2_MPORT_45_data = 1'h0;
  assign ram_2_MPORT_45_addr = 7'h2d;
  assign ram_2_MPORT_45_mask = 1'h1;
  assign ram_2_MPORT_45_en = reset;
  assign ram_2_MPORT_46_data = 1'h0;
  assign ram_2_MPORT_46_addr = 7'h2e;
  assign ram_2_MPORT_46_mask = 1'h1;
  assign ram_2_MPORT_46_en = reset;
  assign ram_2_MPORT_47_data = 1'h0;
  assign ram_2_MPORT_47_addr = 7'h2f;
  assign ram_2_MPORT_47_mask = 1'h1;
  assign ram_2_MPORT_47_en = reset;
  assign ram_2_MPORT_48_data = 1'h0;
  assign ram_2_MPORT_48_addr = 7'h30;
  assign ram_2_MPORT_48_mask = 1'h1;
  assign ram_2_MPORT_48_en = reset;
  assign ram_2_MPORT_49_data = 1'h0;
  assign ram_2_MPORT_49_addr = 7'h31;
  assign ram_2_MPORT_49_mask = 1'h1;
  assign ram_2_MPORT_49_en = reset;
  assign ram_2_MPORT_50_data = 1'h0;
  assign ram_2_MPORT_50_addr = 7'h32;
  assign ram_2_MPORT_50_mask = 1'h1;
  assign ram_2_MPORT_50_en = reset;
  assign ram_2_MPORT_51_data = 1'h0;
  assign ram_2_MPORT_51_addr = 7'h33;
  assign ram_2_MPORT_51_mask = 1'h1;
  assign ram_2_MPORT_51_en = reset;
  assign ram_2_MPORT_52_data = 1'h0;
  assign ram_2_MPORT_52_addr = 7'h34;
  assign ram_2_MPORT_52_mask = 1'h1;
  assign ram_2_MPORT_52_en = reset;
  assign ram_2_MPORT_53_data = 1'h0;
  assign ram_2_MPORT_53_addr = 7'h35;
  assign ram_2_MPORT_53_mask = 1'h1;
  assign ram_2_MPORT_53_en = reset;
  assign ram_2_MPORT_54_data = 1'h0;
  assign ram_2_MPORT_54_addr = 7'h36;
  assign ram_2_MPORT_54_mask = 1'h1;
  assign ram_2_MPORT_54_en = reset;
  assign ram_2_MPORT_55_data = 1'h0;
  assign ram_2_MPORT_55_addr = 7'h37;
  assign ram_2_MPORT_55_mask = 1'h1;
  assign ram_2_MPORT_55_en = reset;
  assign ram_2_MPORT_56_data = 1'h0;
  assign ram_2_MPORT_56_addr = 7'h38;
  assign ram_2_MPORT_56_mask = 1'h1;
  assign ram_2_MPORT_56_en = reset;
  assign ram_2_MPORT_57_data = 1'h0;
  assign ram_2_MPORT_57_addr = 7'h39;
  assign ram_2_MPORT_57_mask = 1'h1;
  assign ram_2_MPORT_57_en = reset;
  assign ram_2_MPORT_58_data = 1'h0;
  assign ram_2_MPORT_58_addr = 7'h3a;
  assign ram_2_MPORT_58_mask = 1'h1;
  assign ram_2_MPORT_58_en = reset;
  assign ram_2_MPORT_59_data = 1'h0;
  assign ram_2_MPORT_59_addr = 7'h3b;
  assign ram_2_MPORT_59_mask = 1'h1;
  assign ram_2_MPORT_59_en = reset;
  assign ram_2_MPORT_60_data = 1'h0;
  assign ram_2_MPORT_60_addr = 7'h3c;
  assign ram_2_MPORT_60_mask = 1'h1;
  assign ram_2_MPORT_60_en = reset;
  assign ram_2_MPORT_61_data = 1'h0;
  assign ram_2_MPORT_61_addr = 7'h3d;
  assign ram_2_MPORT_61_mask = 1'h1;
  assign ram_2_MPORT_61_en = reset;
  assign ram_2_MPORT_62_data = 1'h0;
  assign ram_2_MPORT_62_addr = 7'h3e;
  assign ram_2_MPORT_62_mask = 1'h1;
  assign ram_2_MPORT_62_en = reset;
  assign ram_2_MPORT_63_data = 1'h0;
  assign ram_2_MPORT_63_addr = 7'h3f;
  assign ram_2_MPORT_63_mask = 1'h1;
  assign ram_2_MPORT_63_en = reset;
  assign ram_2_MPORT_64_data = 1'h0;
  assign ram_2_MPORT_64_addr = 7'h40;
  assign ram_2_MPORT_64_mask = 1'h1;
  assign ram_2_MPORT_64_en = reset;
  assign ram_2_MPORT_65_data = 1'h0;
  assign ram_2_MPORT_65_addr = 7'h41;
  assign ram_2_MPORT_65_mask = 1'h1;
  assign ram_2_MPORT_65_en = reset;
  assign ram_2_MPORT_66_data = 1'h0;
  assign ram_2_MPORT_66_addr = 7'h42;
  assign ram_2_MPORT_66_mask = 1'h1;
  assign ram_2_MPORT_66_en = reset;
  assign ram_2_MPORT_67_data = 1'h0;
  assign ram_2_MPORT_67_addr = 7'h43;
  assign ram_2_MPORT_67_mask = 1'h1;
  assign ram_2_MPORT_67_en = reset;
  assign ram_2_MPORT_68_data = 1'h0;
  assign ram_2_MPORT_68_addr = 7'h44;
  assign ram_2_MPORT_68_mask = 1'h1;
  assign ram_2_MPORT_68_en = reset;
  assign ram_2_MPORT_69_data = 1'h0;
  assign ram_2_MPORT_69_addr = 7'h45;
  assign ram_2_MPORT_69_mask = 1'h1;
  assign ram_2_MPORT_69_en = reset;
  assign ram_2_MPORT_70_data = 1'h0;
  assign ram_2_MPORT_70_addr = 7'h46;
  assign ram_2_MPORT_70_mask = 1'h1;
  assign ram_2_MPORT_70_en = reset;
  assign ram_2_MPORT_71_data = 1'h0;
  assign ram_2_MPORT_71_addr = 7'h47;
  assign ram_2_MPORT_71_mask = 1'h1;
  assign ram_2_MPORT_71_en = reset;
  assign ram_2_MPORT_72_data = 1'h0;
  assign ram_2_MPORT_72_addr = 7'h48;
  assign ram_2_MPORT_72_mask = 1'h1;
  assign ram_2_MPORT_72_en = reset;
  assign ram_2_MPORT_73_data = 1'h0;
  assign ram_2_MPORT_73_addr = 7'h49;
  assign ram_2_MPORT_73_mask = 1'h1;
  assign ram_2_MPORT_73_en = reset;
  assign ram_2_MPORT_74_data = 1'h0;
  assign ram_2_MPORT_74_addr = 7'h4a;
  assign ram_2_MPORT_74_mask = 1'h1;
  assign ram_2_MPORT_74_en = reset;
  assign ram_2_MPORT_75_data = 1'h0;
  assign ram_2_MPORT_75_addr = 7'h4b;
  assign ram_2_MPORT_75_mask = 1'h1;
  assign ram_2_MPORT_75_en = reset;
  assign ram_2_MPORT_76_data = 1'h0;
  assign ram_2_MPORT_76_addr = 7'h4c;
  assign ram_2_MPORT_76_mask = 1'h1;
  assign ram_2_MPORT_76_en = reset;
  assign ram_2_MPORT_77_data = 1'h0;
  assign ram_2_MPORT_77_addr = 7'h4d;
  assign ram_2_MPORT_77_mask = 1'h1;
  assign ram_2_MPORT_77_en = reset;
  assign ram_2_MPORT_78_data = 1'h0;
  assign ram_2_MPORT_78_addr = 7'h4e;
  assign ram_2_MPORT_78_mask = 1'h1;
  assign ram_2_MPORT_78_en = reset;
  assign ram_2_MPORT_79_data = 1'h0;
  assign ram_2_MPORT_79_addr = 7'h4f;
  assign ram_2_MPORT_79_mask = 1'h1;
  assign ram_2_MPORT_79_en = reset;
  assign ram_2_MPORT_80_data = 1'h0;
  assign ram_2_MPORT_80_addr = 7'h50;
  assign ram_2_MPORT_80_mask = 1'h1;
  assign ram_2_MPORT_80_en = reset;
  assign ram_2_MPORT_81_data = 1'h0;
  assign ram_2_MPORT_81_addr = 7'h51;
  assign ram_2_MPORT_81_mask = 1'h1;
  assign ram_2_MPORT_81_en = reset;
  assign ram_2_MPORT_82_data = 1'h0;
  assign ram_2_MPORT_82_addr = 7'h52;
  assign ram_2_MPORT_82_mask = 1'h1;
  assign ram_2_MPORT_82_en = reset;
  assign ram_2_MPORT_83_data = 1'h0;
  assign ram_2_MPORT_83_addr = 7'h53;
  assign ram_2_MPORT_83_mask = 1'h1;
  assign ram_2_MPORT_83_en = reset;
  assign ram_2_MPORT_84_data = 1'h0;
  assign ram_2_MPORT_84_addr = 7'h54;
  assign ram_2_MPORT_84_mask = 1'h1;
  assign ram_2_MPORT_84_en = reset;
  assign ram_2_MPORT_85_data = 1'h0;
  assign ram_2_MPORT_85_addr = 7'h55;
  assign ram_2_MPORT_85_mask = 1'h1;
  assign ram_2_MPORT_85_en = reset;
  assign ram_2_MPORT_86_data = 1'h0;
  assign ram_2_MPORT_86_addr = 7'h56;
  assign ram_2_MPORT_86_mask = 1'h1;
  assign ram_2_MPORT_86_en = reset;
  assign ram_2_MPORT_87_data = 1'h0;
  assign ram_2_MPORT_87_addr = 7'h57;
  assign ram_2_MPORT_87_mask = 1'h1;
  assign ram_2_MPORT_87_en = reset;
  assign ram_2_MPORT_88_data = 1'h0;
  assign ram_2_MPORT_88_addr = 7'h58;
  assign ram_2_MPORT_88_mask = 1'h1;
  assign ram_2_MPORT_88_en = reset;
  assign ram_2_MPORT_89_data = 1'h0;
  assign ram_2_MPORT_89_addr = 7'h59;
  assign ram_2_MPORT_89_mask = 1'h1;
  assign ram_2_MPORT_89_en = reset;
  assign ram_2_MPORT_90_data = 1'h0;
  assign ram_2_MPORT_90_addr = 7'h5a;
  assign ram_2_MPORT_90_mask = 1'h1;
  assign ram_2_MPORT_90_en = reset;
  assign ram_2_MPORT_91_data = 1'h0;
  assign ram_2_MPORT_91_addr = 7'h5b;
  assign ram_2_MPORT_91_mask = 1'h1;
  assign ram_2_MPORT_91_en = reset;
  assign ram_2_MPORT_92_data = 1'h0;
  assign ram_2_MPORT_92_addr = 7'h5c;
  assign ram_2_MPORT_92_mask = 1'h1;
  assign ram_2_MPORT_92_en = reset;
  assign ram_2_MPORT_93_data = 1'h0;
  assign ram_2_MPORT_93_addr = 7'h5d;
  assign ram_2_MPORT_93_mask = 1'h1;
  assign ram_2_MPORT_93_en = reset;
  assign ram_2_MPORT_94_data = 1'h0;
  assign ram_2_MPORT_94_addr = 7'h5e;
  assign ram_2_MPORT_94_mask = 1'h1;
  assign ram_2_MPORT_94_en = reset;
  assign ram_2_MPORT_95_data = 1'h0;
  assign ram_2_MPORT_95_addr = 7'h5f;
  assign ram_2_MPORT_95_mask = 1'h1;
  assign ram_2_MPORT_95_en = reset;
  assign ram_2_MPORT_96_data = 1'h0;
  assign ram_2_MPORT_96_addr = 7'h60;
  assign ram_2_MPORT_96_mask = 1'h1;
  assign ram_2_MPORT_96_en = reset;
  assign ram_2_MPORT_97_data = 1'h0;
  assign ram_2_MPORT_97_addr = 7'h61;
  assign ram_2_MPORT_97_mask = 1'h1;
  assign ram_2_MPORT_97_en = reset;
  assign ram_2_MPORT_98_data = 1'h0;
  assign ram_2_MPORT_98_addr = 7'h62;
  assign ram_2_MPORT_98_mask = 1'h1;
  assign ram_2_MPORT_98_en = reset;
  assign ram_2_MPORT_99_data = 1'h0;
  assign ram_2_MPORT_99_addr = 7'h63;
  assign ram_2_MPORT_99_mask = 1'h1;
  assign ram_2_MPORT_99_en = reset;
  assign ram_2_MPORT_100_data = 1'h0;
  assign ram_2_MPORT_100_addr = 7'h64;
  assign ram_2_MPORT_100_mask = 1'h1;
  assign ram_2_MPORT_100_en = reset;
  assign ram_2_MPORT_101_data = 1'h0;
  assign ram_2_MPORT_101_addr = 7'h65;
  assign ram_2_MPORT_101_mask = 1'h1;
  assign ram_2_MPORT_101_en = reset;
  assign ram_2_MPORT_102_data = 1'h0;
  assign ram_2_MPORT_102_addr = 7'h66;
  assign ram_2_MPORT_102_mask = 1'h1;
  assign ram_2_MPORT_102_en = reset;
  assign ram_2_MPORT_103_data = 1'h0;
  assign ram_2_MPORT_103_addr = 7'h67;
  assign ram_2_MPORT_103_mask = 1'h1;
  assign ram_2_MPORT_103_en = reset;
  assign ram_2_MPORT_104_data = 1'h0;
  assign ram_2_MPORT_104_addr = 7'h68;
  assign ram_2_MPORT_104_mask = 1'h1;
  assign ram_2_MPORT_104_en = reset;
  assign ram_2_MPORT_105_data = 1'h0;
  assign ram_2_MPORT_105_addr = 7'h69;
  assign ram_2_MPORT_105_mask = 1'h1;
  assign ram_2_MPORT_105_en = reset;
  assign ram_2_MPORT_106_data = 1'h0;
  assign ram_2_MPORT_106_addr = 7'h6a;
  assign ram_2_MPORT_106_mask = 1'h1;
  assign ram_2_MPORT_106_en = reset;
  assign ram_2_MPORT_107_data = 1'h0;
  assign ram_2_MPORT_107_addr = 7'h6b;
  assign ram_2_MPORT_107_mask = 1'h1;
  assign ram_2_MPORT_107_en = reset;
  assign ram_2_MPORT_108_data = 1'h0;
  assign ram_2_MPORT_108_addr = 7'h6c;
  assign ram_2_MPORT_108_mask = 1'h1;
  assign ram_2_MPORT_108_en = reset;
  assign ram_2_MPORT_109_data = 1'h0;
  assign ram_2_MPORT_109_addr = 7'h6d;
  assign ram_2_MPORT_109_mask = 1'h1;
  assign ram_2_MPORT_109_en = reset;
  assign ram_2_MPORT_110_data = 1'h0;
  assign ram_2_MPORT_110_addr = 7'h6e;
  assign ram_2_MPORT_110_mask = 1'h1;
  assign ram_2_MPORT_110_en = reset;
  assign ram_2_MPORT_111_data = 1'h0;
  assign ram_2_MPORT_111_addr = 7'h6f;
  assign ram_2_MPORT_111_mask = 1'h1;
  assign ram_2_MPORT_111_en = reset;
  assign ram_2_MPORT_112_data = 1'h0;
  assign ram_2_MPORT_112_addr = 7'h70;
  assign ram_2_MPORT_112_mask = 1'h1;
  assign ram_2_MPORT_112_en = reset;
  assign ram_2_MPORT_113_data = 1'h0;
  assign ram_2_MPORT_113_addr = 7'h71;
  assign ram_2_MPORT_113_mask = 1'h1;
  assign ram_2_MPORT_113_en = reset;
  assign ram_2_MPORT_114_data = 1'h0;
  assign ram_2_MPORT_114_addr = 7'h72;
  assign ram_2_MPORT_114_mask = 1'h1;
  assign ram_2_MPORT_114_en = reset;
  assign ram_2_MPORT_115_data = 1'h0;
  assign ram_2_MPORT_115_addr = 7'h73;
  assign ram_2_MPORT_115_mask = 1'h1;
  assign ram_2_MPORT_115_en = reset;
  assign ram_2_MPORT_116_data = 1'h0;
  assign ram_2_MPORT_116_addr = 7'h74;
  assign ram_2_MPORT_116_mask = 1'h1;
  assign ram_2_MPORT_116_en = reset;
  assign ram_2_MPORT_117_data = 1'h0;
  assign ram_2_MPORT_117_addr = 7'h75;
  assign ram_2_MPORT_117_mask = 1'h1;
  assign ram_2_MPORT_117_en = reset;
  assign ram_2_MPORT_118_data = 1'h0;
  assign ram_2_MPORT_118_addr = 7'h76;
  assign ram_2_MPORT_118_mask = 1'h1;
  assign ram_2_MPORT_118_en = reset;
  assign ram_2_MPORT_119_data = 1'h0;
  assign ram_2_MPORT_119_addr = 7'h77;
  assign ram_2_MPORT_119_mask = 1'h1;
  assign ram_2_MPORT_119_en = reset;
  assign ram_2_MPORT_120_data = 1'h0;
  assign ram_2_MPORT_120_addr = 7'h78;
  assign ram_2_MPORT_120_mask = 1'h1;
  assign ram_2_MPORT_120_en = reset;
  assign ram_2_MPORT_121_data = 1'h0;
  assign ram_2_MPORT_121_addr = 7'h79;
  assign ram_2_MPORT_121_mask = 1'h1;
  assign ram_2_MPORT_121_en = reset;
  assign ram_2_MPORT_122_data = 1'h0;
  assign ram_2_MPORT_122_addr = 7'h7a;
  assign ram_2_MPORT_122_mask = 1'h1;
  assign ram_2_MPORT_122_en = reset;
  assign ram_2_MPORT_123_data = 1'h0;
  assign ram_2_MPORT_123_addr = 7'h7b;
  assign ram_2_MPORT_123_mask = 1'h1;
  assign ram_2_MPORT_123_en = reset;
  assign ram_2_MPORT_124_data = 1'h0;
  assign ram_2_MPORT_124_addr = 7'h7c;
  assign ram_2_MPORT_124_mask = 1'h1;
  assign ram_2_MPORT_124_en = reset;
  assign ram_2_MPORT_125_data = 1'h0;
  assign ram_2_MPORT_125_addr = 7'h7d;
  assign ram_2_MPORT_125_mask = 1'h1;
  assign ram_2_MPORT_125_en = reset;
  assign ram_2_MPORT_126_data = 1'h0;
  assign ram_2_MPORT_126_addr = 7'h7e;
  assign ram_2_MPORT_126_mask = 1'h1;
  assign ram_2_MPORT_126_en = reset;
  assign ram_2_MPORT_127_data = 1'h0;
  assign ram_2_MPORT_127_addr = 7'h7f;
  assign ram_2_MPORT_127_mask = 1'h1;
  assign ram_2_MPORT_127_en = reset;
  assign ram_2_MPORT_128_data = 1'h1;
  assign ram_2_MPORT_128_addr = io_addr;
  assign ram_2_MPORT_128_mask = io_wmask[2];
  assign ram_2_MPORT_128_en = io_rw;
  assign ram_3_io_rdata_MPORT_en = ram_3_io_rdata_MPORT_en_pipe_0;
  assign ram_3_io_rdata_MPORT_addr = ram_3_io_rdata_MPORT_addr_pipe_0;
  assign ram_3_io_rdata_MPORT_data = ram_3[ram_3_io_rdata_MPORT_addr]; // @[SRAM.scala 36:26]
  assign ram_3_MPORT_data = 1'h0;
  assign ram_3_MPORT_addr = 7'h0;
  assign ram_3_MPORT_mask = 1'h1;
  assign ram_3_MPORT_en = reset;
  assign ram_3_MPORT_1_data = 1'h0;
  assign ram_3_MPORT_1_addr = 7'h1;
  assign ram_3_MPORT_1_mask = 1'h1;
  assign ram_3_MPORT_1_en = reset;
  assign ram_3_MPORT_2_data = 1'h0;
  assign ram_3_MPORT_2_addr = 7'h2;
  assign ram_3_MPORT_2_mask = 1'h1;
  assign ram_3_MPORT_2_en = reset;
  assign ram_3_MPORT_3_data = 1'h0;
  assign ram_3_MPORT_3_addr = 7'h3;
  assign ram_3_MPORT_3_mask = 1'h1;
  assign ram_3_MPORT_3_en = reset;
  assign ram_3_MPORT_4_data = 1'h0;
  assign ram_3_MPORT_4_addr = 7'h4;
  assign ram_3_MPORT_4_mask = 1'h1;
  assign ram_3_MPORT_4_en = reset;
  assign ram_3_MPORT_5_data = 1'h0;
  assign ram_3_MPORT_5_addr = 7'h5;
  assign ram_3_MPORT_5_mask = 1'h1;
  assign ram_3_MPORT_5_en = reset;
  assign ram_3_MPORT_6_data = 1'h0;
  assign ram_3_MPORT_6_addr = 7'h6;
  assign ram_3_MPORT_6_mask = 1'h1;
  assign ram_3_MPORT_6_en = reset;
  assign ram_3_MPORT_7_data = 1'h0;
  assign ram_3_MPORT_7_addr = 7'h7;
  assign ram_3_MPORT_7_mask = 1'h1;
  assign ram_3_MPORT_7_en = reset;
  assign ram_3_MPORT_8_data = 1'h0;
  assign ram_3_MPORT_8_addr = 7'h8;
  assign ram_3_MPORT_8_mask = 1'h1;
  assign ram_3_MPORT_8_en = reset;
  assign ram_3_MPORT_9_data = 1'h0;
  assign ram_3_MPORT_9_addr = 7'h9;
  assign ram_3_MPORT_9_mask = 1'h1;
  assign ram_3_MPORT_9_en = reset;
  assign ram_3_MPORT_10_data = 1'h0;
  assign ram_3_MPORT_10_addr = 7'ha;
  assign ram_3_MPORT_10_mask = 1'h1;
  assign ram_3_MPORT_10_en = reset;
  assign ram_3_MPORT_11_data = 1'h0;
  assign ram_3_MPORT_11_addr = 7'hb;
  assign ram_3_MPORT_11_mask = 1'h1;
  assign ram_3_MPORT_11_en = reset;
  assign ram_3_MPORT_12_data = 1'h0;
  assign ram_3_MPORT_12_addr = 7'hc;
  assign ram_3_MPORT_12_mask = 1'h1;
  assign ram_3_MPORT_12_en = reset;
  assign ram_3_MPORT_13_data = 1'h0;
  assign ram_3_MPORT_13_addr = 7'hd;
  assign ram_3_MPORT_13_mask = 1'h1;
  assign ram_3_MPORT_13_en = reset;
  assign ram_3_MPORT_14_data = 1'h0;
  assign ram_3_MPORT_14_addr = 7'he;
  assign ram_3_MPORT_14_mask = 1'h1;
  assign ram_3_MPORT_14_en = reset;
  assign ram_3_MPORT_15_data = 1'h0;
  assign ram_3_MPORT_15_addr = 7'hf;
  assign ram_3_MPORT_15_mask = 1'h1;
  assign ram_3_MPORT_15_en = reset;
  assign ram_3_MPORT_16_data = 1'h0;
  assign ram_3_MPORT_16_addr = 7'h10;
  assign ram_3_MPORT_16_mask = 1'h1;
  assign ram_3_MPORT_16_en = reset;
  assign ram_3_MPORT_17_data = 1'h0;
  assign ram_3_MPORT_17_addr = 7'h11;
  assign ram_3_MPORT_17_mask = 1'h1;
  assign ram_3_MPORT_17_en = reset;
  assign ram_3_MPORT_18_data = 1'h0;
  assign ram_3_MPORT_18_addr = 7'h12;
  assign ram_3_MPORT_18_mask = 1'h1;
  assign ram_3_MPORT_18_en = reset;
  assign ram_3_MPORT_19_data = 1'h0;
  assign ram_3_MPORT_19_addr = 7'h13;
  assign ram_3_MPORT_19_mask = 1'h1;
  assign ram_3_MPORT_19_en = reset;
  assign ram_3_MPORT_20_data = 1'h0;
  assign ram_3_MPORT_20_addr = 7'h14;
  assign ram_3_MPORT_20_mask = 1'h1;
  assign ram_3_MPORT_20_en = reset;
  assign ram_3_MPORT_21_data = 1'h0;
  assign ram_3_MPORT_21_addr = 7'h15;
  assign ram_3_MPORT_21_mask = 1'h1;
  assign ram_3_MPORT_21_en = reset;
  assign ram_3_MPORT_22_data = 1'h0;
  assign ram_3_MPORT_22_addr = 7'h16;
  assign ram_3_MPORT_22_mask = 1'h1;
  assign ram_3_MPORT_22_en = reset;
  assign ram_3_MPORT_23_data = 1'h0;
  assign ram_3_MPORT_23_addr = 7'h17;
  assign ram_3_MPORT_23_mask = 1'h1;
  assign ram_3_MPORT_23_en = reset;
  assign ram_3_MPORT_24_data = 1'h0;
  assign ram_3_MPORT_24_addr = 7'h18;
  assign ram_3_MPORT_24_mask = 1'h1;
  assign ram_3_MPORT_24_en = reset;
  assign ram_3_MPORT_25_data = 1'h0;
  assign ram_3_MPORT_25_addr = 7'h19;
  assign ram_3_MPORT_25_mask = 1'h1;
  assign ram_3_MPORT_25_en = reset;
  assign ram_3_MPORT_26_data = 1'h0;
  assign ram_3_MPORT_26_addr = 7'h1a;
  assign ram_3_MPORT_26_mask = 1'h1;
  assign ram_3_MPORT_26_en = reset;
  assign ram_3_MPORT_27_data = 1'h0;
  assign ram_3_MPORT_27_addr = 7'h1b;
  assign ram_3_MPORT_27_mask = 1'h1;
  assign ram_3_MPORT_27_en = reset;
  assign ram_3_MPORT_28_data = 1'h0;
  assign ram_3_MPORT_28_addr = 7'h1c;
  assign ram_3_MPORT_28_mask = 1'h1;
  assign ram_3_MPORT_28_en = reset;
  assign ram_3_MPORT_29_data = 1'h0;
  assign ram_3_MPORT_29_addr = 7'h1d;
  assign ram_3_MPORT_29_mask = 1'h1;
  assign ram_3_MPORT_29_en = reset;
  assign ram_3_MPORT_30_data = 1'h0;
  assign ram_3_MPORT_30_addr = 7'h1e;
  assign ram_3_MPORT_30_mask = 1'h1;
  assign ram_3_MPORT_30_en = reset;
  assign ram_3_MPORT_31_data = 1'h0;
  assign ram_3_MPORT_31_addr = 7'h1f;
  assign ram_3_MPORT_31_mask = 1'h1;
  assign ram_3_MPORT_31_en = reset;
  assign ram_3_MPORT_32_data = 1'h0;
  assign ram_3_MPORT_32_addr = 7'h20;
  assign ram_3_MPORT_32_mask = 1'h1;
  assign ram_3_MPORT_32_en = reset;
  assign ram_3_MPORT_33_data = 1'h0;
  assign ram_3_MPORT_33_addr = 7'h21;
  assign ram_3_MPORT_33_mask = 1'h1;
  assign ram_3_MPORT_33_en = reset;
  assign ram_3_MPORT_34_data = 1'h0;
  assign ram_3_MPORT_34_addr = 7'h22;
  assign ram_3_MPORT_34_mask = 1'h1;
  assign ram_3_MPORT_34_en = reset;
  assign ram_3_MPORT_35_data = 1'h0;
  assign ram_3_MPORT_35_addr = 7'h23;
  assign ram_3_MPORT_35_mask = 1'h1;
  assign ram_3_MPORT_35_en = reset;
  assign ram_3_MPORT_36_data = 1'h0;
  assign ram_3_MPORT_36_addr = 7'h24;
  assign ram_3_MPORT_36_mask = 1'h1;
  assign ram_3_MPORT_36_en = reset;
  assign ram_3_MPORT_37_data = 1'h0;
  assign ram_3_MPORT_37_addr = 7'h25;
  assign ram_3_MPORT_37_mask = 1'h1;
  assign ram_3_MPORT_37_en = reset;
  assign ram_3_MPORT_38_data = 1'h0;
  assign ram_3_MPORT_38_addr = 7'h26;
  assign ram_3_MPORT_38_mask = 1'h1;
  assign ram_3_MPORT_38_en = reset;
  assign ram_3_MPORT_39_data = 1'h0;
  assign ram_3_MPORT_39_addr = 7'h27;
  assign ram_3_MPORT_39_mask = 1'h1;
  assign ram_3_MPORT_39_en = reset;
  assign ram_3_MPORT_40_data = 1'h0;
  assign ram_3_MPORT_40_addr = 7'h28;
  assign ram_3_MPORT_40_mask = 1'h1;
  assign ram_3_MPORT_40_en = reset;
  assign ram_3_MPORT_41_data = 1'h0;
  assign ram_3_MPORT_41_addr = 7'h29;
  assign ram_3_MPORT_41_mask = 1'h1;
  assign ram_3_MPORT_41_en = reset;
  assign ram_3_MPORT_42_data = 1'h0;
  assign ram_3_MPORT_42_addr = 7'h2a;
  assign ram_3_MPORT_42_mask = 1'h1;
  assign ram_3_MPORT_42_en = reset;
  assign ram_3_MPORT_43_data = 1'h0;
  assign ram_3_MPORT_43_addr = 7'h2b;
  assign ram_3_MPORT_43_mask = 1'h1;
  assign ram_3_MPORT_43_en = reset;
  assign ram_3_MPORT_44_data = 1'h0;
  assign ram_3_MPORT_44_addr = 7'h2c;
  assign ram_3_MPORT_44_mask = 1'h1;
  assign ram_3_MPORT_44_en = reset;
  assign ram_3_MPORT_45_data = 1'h0;
  assign ram_3_MPORT_45_addr = 7'h2d;
  assign ram_3_MPORT_45_mask = 1'h1;
  assign ram_3_MPORT_45_en = reset;
  assign ram_3_MPORT_46_data = 1'h0;
  assign ram_3_MPORT_46_addr = 7'h2e;
  assign ram_3_MPORT_46_mask = 1'h1;
  assign ram_3_MPORT_46_en = reset;
  assign ram_3_MPORT_47_data = 1'h0;
  assign ram_3_MPORT_47_addr = 7'h2f;
  assign ram_3_MPORT_47_mask = 1'h1;
  assign ram_3_MPORT_47_en = reset;
  assign ram_3_MPORT_48_data = 1'h0;
  assign ram_3_MPORT_48_addr = 7'h30;
  assign ram_3_MPORT_48_mask = 1'h1;
  assign ram_3_MPORT_48_en = reset;
  assign ram_3_MPORT_49_data = 1'h0;
  assign ram_3_MPORT_49_addr = 7'h31;
  assign ram_3_MPORT_49_mask = 1'h1;
  assign ram_3_MPORT_49_en = reset;
  assign ram_3_MPORT_50_data = 1'h0;
  assign ram_3_MPORT_50_addr = 7'h32;
  assign ram_3_MPORT_50_mask = 1'h1;
  assign ram_3_MPORT_50_en = reset;
  assign ram_3_MPORT_51_data = 1'h0;
  assign ram_3_MPORT_51_addr = 7'h33;
  assign ram_3_MPORT_51_mask = 1'h1;
  assign ram_3_MPORT_51_en = reset;
  assign ram_3_MPORT_52_data = 1'h0;
  assign ram_3_MPORT_52_addr = 7'h34;
  assign ram_3_MPORT_52_mask = 1'h1;
  assign ram_3_MPORT_52_en = reset;
  assign ram_3_MPORT_53_data = 1'h0;
  assign ram_3_MPORT_53_addr = 7'h35;
  assign ram_3_MPORT_53_mask = 1'h1;
  assign ram_3_MPORT_53_en = reset;
  assign ram_3_MPORT_54_data = 1'h0;
  assign ram_3_MPORT_54_addr = 7'h36;
  assign ram_3_MPORT_54_mask = 1'h1;
  assign ram_3_MPORT_54_en = reset;
  assign ram_3_MPORT_55_data = 1'h0;
  assign ram_3_MPORT_55_addr = 7'h37;
  assign ram_3_MPORT_55_mask = 1'h1;
  assign ram_3_MPORT_55_en = reset;
  assign ram_3_MPORT_56_data = 1'h0;
  assign ram_3_MPORT_56_addr = 7'h38;
  assign ram_3_MPORT_56_mask = 1'h1;
  assign ram_3_MPORT_56_en = reset;
  assign ram_3_MPORT_57_data = 1'h0;
  assign ram_3_MPORT_57_addr = 7'h39;
  assign ram_3_MPORT_57_mask = 1'h1;
  assign ram_3_MPORT_57_en = reset;
  assign ram_3_MPORT_58_data = 1'h0;
  assign ram_3_MPORT_58_addr = 7'h3a;
  assign ram_3_MPORT_58_mask = 1'h1;
  assign ram_3_MPORT_58_en = reset;
  assign ram_3_MPORT_59_data = 1'h0;
  assign ram_3_MPORT_59_addr = 7'h3b;
  assign ram_3_MPORT_59_mask = 1'h1;
  assign ram_3_MPORT_59_en = reset;
  assign ram_3_MPORT_60_data = 1'h0;
  assign ram_3_MPORT_60_addr = 7'h3c;
  assign ram_3_MPORT_60_mask = 1'h1;
  assign ram_3_MPORT_60_en = reset;
  assign ram_3_MPORT_61_data = 1'h0;
  assign ram_3_MPORT_61_addr = 7'h3d;
  assign ram_3_MPORT_61_mask = 1'h1;
  assign ram_3_MPORT_61_en = reset;
  assign ram_3_MPORT_62_data = 1'h0;
  assign ram_3_MPORT_62_addr = 7'h3e;
  assign ram_3_MPORT_62_mask = 1'h1;
  assign ram_3_MPORT_62_en = reset;
  assign ram_3_MPORT_63_data = 1'h0;
  assign ram_3_MPORT_63_addr = 7'h3f;
  assign ram_3_MPORT_63_mask = 1'h1;
  assign ram_3_MPORT_63_en = reset;
  assign ram_3_MPORT_64_data = 1'h0;
  assign ram_3_MPORT_64_addr = 7'h40;
  assign ram_3_MPORT_64_mask = 1'h1;
  assign ram_3_MPORT_64_en = reset;
  assign ram_3_MPORT_65_data = 1'h0;
  assign ram_3_MPORT_65_addr = 7'h41;
  assign ram_3_MPORT_65_mask = 1'h1;
  assign ram_3_MPORT_65_en = reset;
  assign ram_3_MPORT_66_data = 1'h0;
  assign ram_3_MPORT_66_addr = 7'h42;
  assign ram_3_MPORT_66_mask = 1'h1;
  assign ram_3_MPORT_66_en = reset;
  assign ram_3_MPORT_67_data = 1'h0;
  assign ram_3_MPORT_67_addr = 7'h43;
  assign ram_3_MPORT_67_mask = 1'h1;
  assign ram_3_MPORT_67_en = reset;
  assign ram_3_MPORT_68_data = 1'h0;
  assign ram_3_MPORT_68_addr = 7'h44;
  assign ram_3_MPORT_68_mask = 1'h1;
  assign ram_3_MPORT_68_en = reset;
  assign ram_3_MPORT_69_data = 1'h0;
  assign ram_3_MPORT_69_addr = 7'h45;
  assign ram_3_MPORT_69_mask = 1'h1;
  assign ram_3_MPORT_69_en = reset;
  assign ram_3_MPORT_70_data = 1'h0;
  assign ram_3_MPORT_70_addr = 7'h46;
  assign ram_3_MPORT_70_mask = 1'h1;
  assign ram_3_MPORT_70_en = reset;
  assign ram_3_MPORT_71_data = 1'h0;
  assign ram_3_MPORT_71_addr = 7'h47;
  assign ram_3_MPORT_71_mask = 1'h1;
  assign ram_3_MPORT_71_en = reset;
  assign ram_3_MPORT_72_data = 1'h0;
  assign ram_3_MPORT_72_addr = 7'h48;
  assign ram_3_MPORT_72_mask = 1'h1;
  assign ram_3_MPORT_72_en = reset;
  assign ram_3_MPORT_73_data = 1'h0;
  assign ram_3_MPORT_73_addr = 7'h49;
  assign ram_3_MPORT_73_mask = 1'h1;
  assign ram_3_MPORT_73_en = reset;
  assign ram_3_MPORT_74_data = 1'h0;
  assign ram_3_MPORT_74_addr = 7'h4a;
  assign ram_3_MPORT_74_mask = 1'h1;
  assign ram_3_MPORT_74_en = reset;
  assign ram_3_MPORT_75_data = 1'h0;
  assign ram_3_MPORT_75_addr = 7'h4b;
  assign ram_3_MPORT_75_mask = 1'h1;
  assign ram_3_MPORT_75_en = reset;
  assign ram_3_MPORT_76_data = 1'h0;
  assign ram_3_MPORT_76_addr = 7'h4c;
  assign ram_3_MPORT_76_mask = 1'h1;
  assign ram_3_MPORT_76_en = reset;
  assign ram_3_MPORT_77_data = 1'h0;
  assign ram_3_MPORT_77_addr = 7'h4d;
  assign ram_3_MPORT_77_mask = 1'h1;
  assign ram_3_MPORT_77_en = reset;
  assign ram_3_MPORT_78_data = 1'h0;
  assign ram_3_MPORT_78_addr = 7'h4e;
  assign ram_3_MPORT_78_mask = 1'h1;
  assign ram_3_MPORT_78_en = reset;
  assign ram_3_MPORT_79_data = 1'h0;
  assign ram_3_MPORT_79_addr = 7'h4f;
  assign ram_3_MPORT_79_mask = 1'h1;
  assign ram_3_MPORT_79_en = reset;
  assign ram_3_MPORT_80_data = 1'h0;
  assign ram_3_MPORT_80_addr = 7'h50;
  assign ram_3_MPORT_80_mask = 1'h1;
  assign ram_3_MPORT_80_en = reset;
  assign ram_3_MPORT_81_data = 1'h0;
  assign ram_3_MPORT_81_addr = 7'h51;
  assign ram_3_MPORT_81_mask = 1'h1;
  assign ram_3_MPORT_81_en = reset;
  assign ram_3_MPORT_82_data = 1'h0;
  assign ram_3_MPORT_82_addr = 7'h52;
  assign ram_3_MPORT_82_mask = 1'h1;
  assign ram_3_MPORT_82_en = reset;
  assign ram_3_MPORT_83_data = 1'h0;
  assign ram_3_MPORT_83_addr = 7'h53;
  assign ram_3_MPORT_83_mask = 1'h1;
  assign ram_3_MPORT_83_en = reset;
  assign ram_3_MPORT_84_data = 1'h0;
  assign ram_3_MPORT_84_addr = 7'h54;
  assign ram_3_MPORT_84_mask = 1'h1;
  assign ram_3_MPORT_84_en = reset;
  assign ram_3_MPORT_85_data = 1'h0;
  assign ram_3_MPORT_85_addr = 7'h55;
  assign ram_3_MPORT_85_mask = 1'h1;
  assign ram_3_MPORT_85_en = reset;
  assign ram_3_MPORT_86_data = 1'h0;
  assign ram_3_MPORT_86_addr = 7'h56;
  assign ram_3_MPORT_86_mask = 1'h1;
  assign ram_3_MPORT_86_en = reset;
  assign ram_3_MPORT_87_data = 1'h0;
  assign ram_3_MPORT_87_addr = 7'h57;
  assign ram_3_MPORT_87_mask = 1'h1;
  assign ram_3_MPORT_87_en = reset;
  assign ram_3_MPORT_88_data = 1'h0;
  assign ram_3_MPORT_88_addr = 7'h58;
  assign ram_3_MPORT_88_mask = 1'h1;
  assign ram_3_MPORT_88_en = reset;
  assign ram_3_MPORT_89_data = 1'h0;
  assign ram_3_MPORT_89_addr = 7'h59;
  assign ram_3_MPORT_89_mask = 1'h1;
  assign ram_3_MPORT_89_en = reset;
  assign ram_3_MPORT_90_data = 1'h0;
  assign ram_3_MPORT_90_addr = 7'h5a;
  assign ram_3_MPORT_90_mask = 1'h1;
  assign ram_3_MPORT_90_en = reset;
  assign ram_3_MPORT_91_data = 1'h0;
  assign ram_3_MPORT_91_addr = 7'h5b;
  assign ram_3_MPORT_91_mask = 1'h1;
  assign ram_3_MPORT_91_en = reset;
  assign ram_3_MPORT_92_data = 1'h0;
  assign ram_3_MPORT_92_addr = 7'h5c;
  assign ram_3_MPORT_92_mask = 1'h1;
  assign ram_3_MPORT_92_en = reset;
  assign ram_3_MPORT_93_data = 1'h0;
  assign ram_3_MPORT_93_addr = 7'h5d;
  assign ram_3_MPORT_93_mask = 1'h1;
  assign ram_3_MPORT_93_en = reset;
  assign ram_3_MPORT_94_data = 1'h0;
  assign ram_3_MPORT_94_addr = 7'h5e;
  assign ram_3_MPORT_94_mask = 1'h1;
  assign ram_3_MPORT_94_en = reset;
  assign ram_3_MPORT_95_data = 1'h0;
  assign ram_3_MPORT_95_addr = 7'h5f;
  assign ram_3_MPORT_95_mask = 1'h1;
  assign ram_3_MPORT_95_en = reset;
  assign ram_3_MPORT_96_data = 1'h0;
  assign ram_3_MPORT_96_addr = 7'h60;
  assign ram_3_MPORT_96_mask = 1'h1;
  assign ram_3_MPORT_96_en = reset;
  assign ram_3_MPORT_97_data = 1'h0;
  assign ram_3_MPORT_97_addr = 7'h61;
  assign ram_3_MPORT_97_mask = 1'h1;
  assign ram_3_MPORT_97_en = reset;
  assign ram_3_MPORT_98_data = 1'h0;
  assign ram_3_MPORT_98_addr = 7'h62;
  assign ram_3_MPORT_98_mask = 1'h1;
  assign ram_3_MPORT_98_en = reset;
  assign ram_3_MPORT_99_data = 1'h0;
  assign ram_3_MPORT_99_addr = 7'h63;
  assign ram_3_MPORT_99_mask = 1'h1;
  assign ram_3_MPORT_99_en = reset;
  assign ram_3_MPORT_100_data = 1'h0;
  assign ram_3_MPORT_100_addr = 7'h64;
  assign ram_3_MPORT_100_mask = 1'h1;
  assign ram_3_MPORT_100_en = reset;
  assign ram_3_MPORT_101_data = 1'h0;
  assign ram_3_MPORT_101_addr = 7'h65;
  assign ram_3_MPORT_101_mask = 1'h1;
  assign ram_3_MPORT_101_en = reset;
  assign ram_3_MPORT_102_data = 1'h0;
  assign ram_3_MPORT_102_addr = 7'h66;
  assign ram_3_MPORT_102_mask = 1'h1;
  assign ram_3_MPORT_102_en = reset;
  assign ram_3_MPORT_103_data = 1'h0;
  assign ram_3_MPORT_103_addr = 7'h67;
  assign ram_3_MPORT_103_mask = 1'h1;
  assign ram_3_MPORT_103_en = reset;
  assign ram_3_MPORT_104_data = 1'h0;
  assign ram_3_MPORT_104_addr = 7'h68;
  assign ram_3_MPORT_104_mask = 1'h1;
  assign ram_3_MPORT_104_en = reset;
  assign ram_3_MPORT_105_data = 1'h0;
  assign ram_3_MPORT_105_addr = 7'h69;
  assign ram_3_MPORT_105_mask = 1'h1;
  assign ram_3_MPORT_105_en = reset;
  assign ram_3_MPORT_106_data = 1'h0;
  assign ram_3_MPORT_106_addr = 7'h6a;
  assign ram_3_MPORT_106_mask = 1'h1;
  assign ram_3_MPORT_106_en = reset;
  assign ram_3_MPORT_107_data = 1'h0;
  assign ram_3_MPORT_107_addr = 7'h6b;
  assign ram_3_MPORT_107_mask = 1'h1;
  assign ram_3_MPORT_107_en = reset;
  assign ram_3_MPORT_108_data = 1'h0;
  assign ram_3_MPORT_108_addr = 7'h6c;
  assign ram_3_MPORT_108_mask = 1'h1;
  assign ram_3_MPORT_108_en = reset;
  assign ram_3_MPORT_109_data = 1'h0;
  assign ram_3_MPORT_109_addr = 7'h6d;
  assign ram_3_MPORT_109_mask = 1'h1;
  assign ram_3_MPORT_109_en = reset;
  assign ram_3_MPORT_110_data = 1'h0;
  assign ram_3_MPORT_110_addr = 7'h6e;
  assign ram_3_MPORT_110_mask = 1'h1;
  assign ram_3_MPORT_110_en = reset;
  assign ram_3_MPORT_111_data = 1'h0;
  assign ram_3_MPORT_111_addr = 7'h6f;
  assign ram_3_MPORT_111_mask = 1'h1;
  assign ram_3_MPORT_111_en = reset;
  assign ram_3_MPORT_112_data = 1'h0;
  assign ram_3_MPORT_112_addr = 7'h70;
  assign ram_3_MPORT_112_mask = 1'h1;
  assign ram_3_MPORT_112_en = reset;
  assign ram_3_MPORT_113_data = 1'h0;
  assign ram_3_MPORT_113_addr = 7'h71;
  assign ram_3_MPORT_113_mask = 1'h1;
  assign ram_3_MPORT_113_en = reset;
  assign ram_3_MPORT_114_data = 1'h0;
  assign ram_3_MPORT_114_addr = 7'h72;
  assign ram_3_MPORT_114_mask = 1'h1;
  assign ram_3_MPORT_114_en = reset;
  assign ram_3_MPORT_115_data = 1'h0;
  assign ram_3_MPORT_115_addr = 7'h73;
  assign ram_3_MPORT_115_mask = 1'h1;
  assign ram_3_MPORT_115_en = reset;
  assign ram_3_MPORT_116_data = 1'h0;
  assign ram_3_MPORT_116_addr = 7'h74;
  assign ram_3_MPORT_116_mask = 1'h1;
  assign ram_3_MPORT_116_en = reset;
  assign ram_3_MPORT_117_data = 1'h0;
  assign ram_3_MPORT_117_addr = 7'h75;
  assign ram_3_MPORT_117_mask = 1'h1;
  assign ram_3_MPORT_117_en = reset;
  assign ram_3_MPORT_118_data = 1'h0;
  assign ram_3_MPORT_118_addr = 7'h76;
  assign ram_3_MPORT_118_mask = 1'h1;
  assign ram_3_MPORT_118_en = reset;
  assign ram_3_MPORT_119_data = 1'h0;
  assign ram_3_MPORT_119_addr = 7'h77;
  assign ram_3_MPORT_119_mask = 1'h1;
  assign ram_3_MPORT_119_en = reset;
  assign ram_3_MPORT_120_data = 1'h0;
  assign ram_3_MPORT_120_addr = 7'h78;
  assign ram_3_MPORT_120_mask = 1'h1;
  assign ram_3_MPORT_120_en = reset;
  assign ram_3_MPORT_121_data = 1'h0;
  assign ram_3_MPORT_121_addr = 7'h79;
  assign ram_3_MPORT_121_mask = 1'h1;
  assign ram_3_MPORT_121_en = reset;
  assign ram_3_MPORT_122_data = 1'h0;
  assign ram_3_MPORT_122_addr = 7'h7a;
  assign ram_3_MPORT_122_mask = 1'h1;
  assign ram_3_MPORT_122_en = reset;
  assign ram_3_MPORT_123_data = 1'h0;
  assign ram_3_MPORT_123_addr = 7'h7b;
  assign ram_3_MPORT_123_mask = 1'h1;
  assign ram_3_MPORT_123_en = reset;
  assign ram_3_MPORT_124_data = 1'h0;
  assign ram_3_MPORT_124_addr = 7'h7c;
  assign ram_3_MPORT_124_mask = 1'h1;
  assign ram_3_MPORT_124_en = reset;
  assign ram_3_MPORT_125_data = 1'h0;
  assign ram_3_MPORT_125_addr = 7'h7d;
  assign ram_3_MPORT_125_mask = 1'h1;
  assign ram_3_MPORT_125_en = reset;
  assign ram_3_MPORT_126_data = 1'h0;
  assign ram_3_MPORT_126_addr = 7'h7e;
  assign ram_3_MPORT_126_mask = 1'h1;
  assign ram_3_MPORT_126_en = reset;
  assign ram_3_MPORT_127_data = 1'h0;
  assign ram_3_MPORT_127_addr = 7'h7f;
  assign ram_3_MPORT_127_mask = 1'h1;
  assign ram_3_MPORT_127_en = reset;
  assign ram_3_MPORT_128_data = 1'h1;
  assign ram_3_MPORT_128_addr = io_addr;
  assign ram_3_MPORT_128_mask = io_wmask[3];
  assign ram_3_MPORT_128_en = io_rw;
  assign io_rdata = {io_rdata_hi,io_rdata_lo}; // @[SRAM.scala 75:39]
  always @(posedge clock) begin
    if (ram_0_MPORT_en & ram_0_MPORT_mask) begin
      ram_0[ram_0_MPORT_addr] <= ram_0_MPORT_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_1_en & ram_0_MPORT_1_mask) begin
      ram_0[ram_0_MPORT_1_addr] <= ram_0_MPORT_1_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_2_en & ram_0_MPORT_2_mask) begin
      ram_0[ram_0_MPORT_2_addr] <= ram_0_MPORT_2_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_3_en & ram_0_MPORT_3_mask) begin
      ram_0[ram_0_MPORT_3_addr] <= ram_0_MPORT_3_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_4_en & ram_0_MPORT_4_mask) begin
      ram_0[ram_0_MPORT_4_addr] <= ram_0_MPORT_4_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_5_en & ram_0_MPORT_5_mask) begin
      ram_0[ram_0_MPORT_5_addr] <= ram_0_MPORT_5_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_6_en & ram_0_MPORT_6_mask) begin
      ram_0[ram_0_MPORT_6_addr] <= ram_0_MPORT_6_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_7_en & ram_0_MPORT_7_mask) begin
      ram_0[ram_0_MPORT_7_addr] <= ram_0_MPORT_7_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_8_en & ram_0_MPORT_8_mask) begin
      ram_0[ram_0_MPORT_8_addr] <= ram_0_MPORT_8_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_9_en & ram_0_MPORT_9_mask) begin
      ram_0[ram_0_MPORT_9_addr] <= ram_0_MPORT_9_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_10_en & ram_0_MPORT_10_mask) begin
      ram_0[ram_0_MPORT_10_addr] <= ram_0_MPORT_10_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_11_en & ram_0_MPORT_11_mask) begin
      ram_0[ram_0_MPORT_11_addr] <= ram_0_MPORT_11_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_12_en & ram_0_MPORT_12_mask) begin
      ram_0[ram_0_MPORT_12_addr] <= ram_0_MPORT_12_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_13_en & ram_0_MPORT_13_mask) begin
      ram_0[ram_0_MPORT_13_addr] <= ram_0_MPORT_13_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_14_en & ram_0_MPORT_14_mask) begin
      ram_0[ram_0_MPORT_14_addr] <= ram_0_MPORT_14_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_15_en & ram_0_MPORT_15_mask) begin
      ram_0[ram_0_MPORT_15_addr] <= ram_0_MPORT_15_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_16_en & ram_0_MPORT_16_mask) begin
      ram_0[ram_0_MPORT_16_addr] <= ram_0_MPORT_16_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_17_en & ram_0_MPORT_17_mask) begin
      ram_0[ram_0_MPORT_17_addr] <= ram_0_MPORT_17_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_18_en & ram_0_MPORT_18_mask) begin
      ram_0[ram_0_MPORT_18_addr] <= ram_0_MPORT_18_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_19_en & ram_0_MPORT_19_mask) begin
      ram_0[ram_0_MPORT_19_addr] <= ram_0_MPORT_19_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_20_en & ram_0_MPORT_20_mask) begin
      ram_0[ram_0_MPORT_20_addr] <= ram_0_MPORT_20_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_21_en & ram_0_MPORT_21_mask) begin
      ram_0[ram_0_MPORT_21_addr] <= ram_0_MPORT_21_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_22_en & ram_0_MPORT_22_mask) begin
      ram_0[ram_0_MPORT_22_addr] <= ram_0_MPORT_22_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_23_en & ram_0_MPORT_23_mask) begin
      ram_0[ram_0_MPORT_23_addr] <= ram_0_MPORT_23_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_24_en & ram_0_MPORT_24_mask) begin
      ram_0[ram_0_MPORT_24_addr] <= ram_0_MPORT_24_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_25_en & ram_0_MPORT_25_mask) begin
      ram_0[ram_0_MPORT_25_addr] <= ram_0_MPORT_25_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_26_en & ram_0_MPORT_26_mask) begin
      ram_0[ram_0_MPORT_26_addr] <= ram_0_MPORT_26_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_27_en & ram_0_MPORT_27_mask) begin
      ram_0[ram_0_MPORT_27_addr] <= ram_0_MPORT_27_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_28_en & ram_0_MPORT_28_mask) begin
      ram_0[ram_0_MPORT_28_addr] <= ram_0_MPORT_28_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_29_en & ram_0_MPORT_29_mask) begin
      ram_0[ram_0_MPORT_29_addr] <= ram_0_MPORT_29_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_30_en & ram_0_MPORT_30_mask) begin
      ram_0[ram_0_MPORT_30_addr] <= ram_0_MPORT_30_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_31_en & ram_0_MPORT_31_mask) begin
      ram_0[ram_0_MPORT_31_addr] <= ram_0_MPORT_31_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_32_en & ram_0_MPORT_32_mask) begin
      ram_0[ram_0_MPORT_32_addr] <= ram_0_MPORT_32_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_33_en & ram_0_MPORT_33_mask) begin
      ram_0[ram_0_MPORT_33_addr] <= ram_0_MPORT_33_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_34_en & ram_0_MPORT_34_mask) begin
      ram_0[ram_0_MPORT_34_addr] <= ram_0_MPORT_34_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_35_en & ram_0_MPORT_35_mask) begin
      ram_0[ram_0_MPORT_35_addr] <= ram_0_MPORT_35_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_36_en & ram_0_MPORT_36_mask) begin
      ram_0[ram_0_MPORT_36_addr] <= ram_0_MPORT_36_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_37_en & ram_0_MPORT_37_mask) begin
      ram_0[ram_0_MPORT_37_addr] <= ram_0_MPORT_37_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_38_en & ram_0_MPORT_38_mask) begin
      ram_0[ram_0_MPORT_38_addr] <= ram_0_MPORT_38_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_39_en & ram_0_MPORT_39_mask) begin
      ram_0[ram_0_MPORT_39_addr] <= ram_0_MPORT_39_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_40_en & ram_0_MPORT_40_mask) begin
      ram_0[ram_0_MPORT_40_addr] <= ram_0_MPORT_40_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_41_en & ram_0_MPORT_41_mask) begin
      ram_0[ram_0_MPORT_41_addr] <= ram_0_MPORT_41_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_42_en & ram_0_MPORT_42_mask) begin
      ram_0[ram_0_MPORT_42_addr] <= ram_0_MPORT_42_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_43_en & ram_0_MPORT_43_mask) begin
      ram_0[ram_0_MPORT_43_addr] <= ram_0_MPORT_43_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_44_en & ram_0_MPORT_44_mask) begin
      ram_0[ram_0_MPORT_44_addr] <= ram_0_MPORT_44_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_45_en & ram_0_MPORT_45_mask) begin
      ram_0[ram_0_MPORT_45_addr] <= ram_0_MPORT_45_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_46_en & ram_0_MPORT_46_mask) begin
      ram_0[ram_0_MPORT_46_addr] <= ram_0_MPORT_46_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_47_en & ram_0_MPORT_47_mask) begin
      ram_0[ram_0_MPORT_47_addr] <= ram_0_MPORT_47_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_48_en & ram_0_MPORT_48_mask) begin
      ram_0[ram_0_MPORT_48_addr] <= ram_0_MPORT_48_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_49_en & ram_0_MPORT_49_mask) begin
      ram_0[ram_0_MPORT_49_addr] <= ram_0_MPORT_49_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_50_en & ram_0_MPORT_50_mask) begin
      ram_0[ram_0_MPORT_50_addr] <= ram_0_MPORT_50_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_51_en & ram_0_MPORT_51_mask) begin
      ram_0[ram_0_MPORT_51_addr] <= ram_0_MPORT_51_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_52_en & ram_0_MPORT_52_mask) begin
      ram_0[ram_0_MPORT_52_addr] <= ram_0_MPORT_52_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_53_en & ram_0_MPORT_53_mask) begin
      ram_0[ram_0_MPORT_53_addr] <= ram_0_MPORT_53_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_54_en & ram_0_MPORT_54_mask) begin
      ram_0[ram_0_MPORT_54_addr] <= ram_0_MPORT_54_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_55_en & ram_0_MPORT_55_mask) begin
      ram_0[ram_0_MPORT_55_addr] <= ram_0_MPORT_55_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_56_en & ram_0_MPORT_56_mask) begin
      ram_0[ram_0_MPORT_56_addr] <= ram_0_MPORT_56_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_57_en & ram_0_MPORT_57_mask) begin
      ram_0[ram_0_MPORT_57_addr] <= ram_0_MPORT_57_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_58_en & ram_0_MPORT_58_mask) begin
      ram_0[ram_0_MPORT_58_addr] <= ram_0_MPORT_58_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_59_en & ram_0_MPORT_59_mask) begin
      ram_0[ram_0_MPORT_59_addr] <= ram_0_MPORT_59_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_60_en & ram_0_MPORT_60_mask) begin
      ram_0[ram_0_MPORT_60_addr] <= ram_0_MPORT_60_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_61_en & ram_0_MPORT_61_mask) begin
      ram_0[ram_0_MPORT_61_addr] <= ram_0_MPORT_61_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_62_en & ram_0_MPORT_62_mask) begin
      ram_0[ram_0_MPORT_62_addr] <= ram_0_MPORT_62_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_63_en & ram_0_MPORT_63_mask) begin
      ram_0[ram_0_MPORT_63_addr] <= ram_0_MPORT_63_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_64_en & ram_0_MPORT_64_mask) begin
      ram_0[ram_0_MPORT_64_addr] <= ram_0_MPORT_64_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_65_en & ram_0_MPORT_65_mask) begin
      ram_0[ram_0_MPORT_65_addr] <= ram_0_MPORT_65_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_66_en & ram_0_MPORT_66_mask) begin
      ram_0[ram_0_MPORT_66_addr] <= ram_0_MPORT_66_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_67_en & ram_0_MPORT_67_mask) begin
      ram_0[ram_0_MPORT_67_addr] <= ram_0_MPORT_67_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_68_en & ram_0_MPORT_68_mask) begin
      ram_0[ram_0_MPORT_68_addr] <= ram_0_MPORT_68_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_69_en & ram_0_MPORT_69_mask) begin
      ram_0[ram_0_MPORT_69_addr] <= ram_0_MPORT_69_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_70_en & ram_0_MPORT_70_mask) begin
      ram_0[ram_0_MPORT_70_addr] <= ram_0_MPORT_70_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_71_en & ram_0_MPORT_71_mask) begin
      ram_0[ram_0_MPORT_71_addr] <= ram_0_MPORT_71_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_72_en & ram_0_MPORT_72_mask) begin
      ram_0[ram_0_MPORT_72_addr] <= ram_0_MPORT_72_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_73_en & ram_0_MPORT_73_mask) begin
      ram_0[ram_0_MPORT_73_addr] <= ram_0_MPORT_73_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_74_en & ram_0_MPORT_74_mask) begin
      ram_0[ram_0_MPORT_74_addr] <= ram_0_MPORT_74_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_75_en & ram_0_MPORT_75_mask) begin
      ram_0[ram_0_MPORT_75_addr] <= ram_0_MPORT_75_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_76_en & ram_0_MPORT_76_mask) begin
      ram_0[ram_0_MPORT_76_addr] <= ram_0_MPORT_76_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_77_en & ram_0_MPORT_77_mask) begin
      ram_0[ram_0_MPORT_77_addr] <= ram_0_MPORT_77_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_78_en & ram_0_MPORT_78_mask) begin
      ram_0[ram_0_MPORT_78_addr] <= ram_0_MPORT_78_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_79_en & ram_0_MPORT_79_mask) begin
      ram_0[ram_0_MPORT_79_addr] <= ram_0_MPORT_79_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_80_en & ram_0_MPORT_80_mask) begin
      ram_0[ram_0_MPORT_80_addr] <= ram_0_MPORT_80_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_81_en & ram_0_MPORT_81_mask) begin
      ram_0[ram_0_MPORT_81_addr] <= ram_0_MPORT_81_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_82_en & ram_0_MPORT_82_mask) begin
      ram_0[ram_0_MPORT_82_addr] <= ram_0_MPORT_82_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_83_en & ram_0_MPORT_83_mask) begin
      ram_0[ram_0_MPORT_83_addr] <= ram_0_MPORT_83_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_84_en & ram_0_MPORT_84_mask) begin
      ram_0[ram_0_MPORT_84_addr] <= ram_0_MPORT_84_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_85_en & ram_0_MPORT_85_mask) begin
      ram_0[ram_0_MPORT_85_addr] <= ram_0_MPORT_85_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_86_en & ram_0_MPORT_86_mask) begin
      ram_0[ram_0_MPORT_86_addr] <= ram_0_MPORT_86_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_87_en & ram_0_MPORT_87_mask) begin
      ram_0[ram_0_MPORT_87_addr] <= ram_0_MPORT_87_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_88_en & ram_0_MPORT_88_mask) begin
      ram_0[ram_0_MPORT_88_addr] <= ram_0_MPORT_88_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_89_en & ram_0_MPORT_89_mask) begin
      ram_0[ram_0_MPORT_89_addr] <= ram_0_MPORT_89_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_90_en & ram_0_MPORT_90_mask) begin
      ram_0[ram_0_MPORT_90_addr] <= ram_0_MPORT_90_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_91_en & ram_0_MPORT_91_mask) begin
      ram_0[ram_0_MPORT_91_addr] <= ram_0_MPORT_91_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_92_en & ram_0_MPORT_92_mask) begin
      ram_0[ram_0_MPORT_92_addr] <= ram_0_MPORT_92_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_93_en & ram_0_MPORT_93_mask) begin
      ram_0[ram_0_MPORT_93_addr] <= ram_0_MPORT_93_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_94_en & ram_0_MPORT_94_mask) begin
      ram_0[ram_0_MPORT_94_addr] <= ram_0_MPORT_94_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_95_en & ram_0_MPORT_95_mask) begin
      ram_0[ram_0_MPORT_95_addr] <= ram_0_MPORT_95_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_96_en & ram_0_MPORT_96_mask) begin
      ram_0[ram_0_MPORT_96_addr] <= ram_0_MPORT_96_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_97_en & ram_0_MPORT_97_mask) begin
      ram_0[ram_0_MPORT_97_addr] <= ram_0_MPORT_97_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_98_en & ram_0_MPORT_98_mask) begin
      ram_0[ram_0_MPORT_98_addr] <= ram_0_MPORT_98_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_99_en & ram_0_MPORT_99_mask) begin
      ram_0[ram_0_MPORT_99_addr] <= ram_0_MPORT_99_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_100_en & ram_0_MPORT_100_mask) begin
      ram_0[ram_0_MPORT_100_addr] <= ram_0_MPORT_100_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_101_en & ram_0_MPORT_101_mask) begin
      ram_0[ram_0_MPORT_101_addr] <= ram_0_MPORT_101_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_102_en & ram_0_MPORT_102_mask) begin
      ram_0[ram_0_MPORT_102_addr] <= ram_0_MPORT_102_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_103_en & ram_0_MPORT_103_mask) begin
      ram_0[ram_0_MPORT_103_addr] <= ram_0_MPORT_103_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_104_en & ram_0_MPORT_104_mask) begin
      ram_0[ram_0_MPORT_104_addr] <= ram_0_MPORT_104_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_105_en & ram_0_MPORT_105_mask) begin
      ram_0[ram_0_MPORT_105_addr] <= ram_0_MPORT_105_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_106_en & ram_0_MPORT_106_mask) begin
      ram_0[ram_0_MPORT_106_addr] <= ram_0_MPORT_106_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_107_en & ram_0_MPORT_107_mask) begin
      ram_0[ram_0_MPORT_107_addr] <= ram_0_MPORT_107_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_108_en & ram_0_MPORT_108_mask) begin
      ram_0[ram_0_MPORT_108_addr] <= ram_0_MPORT_108_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_109_en & ram_0_MPORT_109_mask) begin
      ram_0[ram_0_MPORT_109_addr] <= ram_0_MPORT_109_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_110_en & ram_0_MPORT_110_mask) begin
      ram_0[ram_0_MPORT_110_addr] <= ram_0_MPORT_110_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_111_en & ram_0_MPORT_111_mask) begin
      ram_0[ram_0_MPORT_111_addr] <= ram_0_MPORT_111_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_112_en & ram_0_MPORT_112_mask) begin
      ram_0[ram_0_MPORT_112_addr] <= ram_0_MPORT_112_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_113_en & ram_0_MPORT_113_mask) begin
      ram_0[ram_0_MPORT_113_addr] <= ram_0_MPORT_113_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_114_en & ram_0_MPORT_114_mask) begin
      ram_0[ram_0_MPORT_114_addr] <= ram_0_MPORT_114_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_115_en & ram_0_MPORT_115_mask) begin
      ram_0[ram_0_MPORT_115_addr] <= ram_0_MPORT_115_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_116_en & ram_0_MPORT_116_mask) begin
      ram_0[ram_0_MPORT_116_addr] <= ram_0_MPORT_116_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_117_en & ram_0_MPORT_117_mask) begin
      ram_0[ram_0_MPORT_117_addr] <= ram_0_MPORT_117_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_118_en & ram_0_MPORT_118_mask) begin
      ram_0[ram_0_MPORT_118_addr] <= ram_0_MPORT_118_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_119_en & ram_0_MPORT_119_mask) begin
      ram_0[ram_0_MPORT_119_addr] <= ram_0_MPORT_119_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_120_en & ram_0_MPORT_120_mask) begin
      ram_0[ram_0_MPORT_120_addr] <= ram_0_MPORT_120_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_121_en & ram_0_MPORT_121_mask) begin
      ram_0[ram_0_MPORT_121_addr] <= ram_0_MPORT_121_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_122_en & ram_0_MPORT_122_mask) begin
      ram_0[ram_0_MPORT_122_addr] <= ram_0_MPORT_122_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_123_en & ram_0_MPORT_123_mask) begin
      ram_0[ram_0_MPORT_123_addr] <= ram_0_MPORT_123_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_124_en & ram_0_MPORT_124_mask) begin
      ram_0[ram_0_MPORT_124_addr] <= ram_0_MPORT_124_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_125_en & ram_0_MPORT_125_mask) begin
      ram_0[ram_0_MPORT_125_addr] <= ram_0_MPORT_125_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_126_en & ram_0_MPORT_126_mask) begin
      ram_0[ram_0_MPORT_126_addr] <= ram_0_MPORT_126_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_127_en & ram_0_MPORT_127_mask) begin
      ram_0[ram_0_MPORT_127_addr] <= ram_0_MPORT_127_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_128_en & ram_0_MPORT_128_mask) begin
      ram_0[ram_0_MPORT_128_addr] <= ram_0_MPORT_128_data; // @[SRAM.scala 36:26]
    end
    if (io_rw) begin
      ram_0_io_rdata_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      ram_0_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    end
    if (io_rw ? 1'h0 : 1'h1) begin
      ram_0_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
    if (ram_1_MPORT_en & ram_1_MPORT_mask) begin
      ram_1[ram_1_MPORT_addr] <= ram_1_MPORT_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_1_en & ram_1_MPORT_1_mask) begin
      ram_1[ram_1_MPORT_1_addr] <= ram_1_MPORT_1_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_2_en & ram_1_MPORT_2_mask) begin
      ram_1[ram_1_MPORT_2_addr] <= ram_1_MPORT_2_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_3_en & ram_1_MPORT_3_mask) begin
      ram_1[ram_1_MPORT_3_addr] <= ram_1_MPORT_3_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_4_en & ram_1_MPORT_4_mask) begin
      ram_1[ram_1_MPORT_4_addr] <= ram_1_MPORT_4_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_5_en & ram_1_MPORT_5_mask) begin
      ram_1[ram_1_MPORT_5_addr] <= ram_1_MPORT_5_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_6_en & ram_1_MPORT_6_mask) begin
      ram_1[ram_1_MPORT_6_addr] <= ram_1_MPORT_6_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_7_en & ram_1_MPORT_7_mask) begin
      ram_1[ram_1_MPORT_7_addr] <= ram_1_MPORT_7_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_8_en & ram_1_MPORT_8_mask) begin
      ram_1[ram_1_MPORT_8_addr] <= ram_1_MPORT_8_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_9_en & ram_1_MPORT_9_mask) begin
      ram_1[ram_1_MPORT_9_addr] <= ram_1_MPORT_9_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_10_en & ram_1_MPORT_10_mask) begin
      ram_1[ram_1_MPORT_10_addr] <= ram_1_MPORT_10_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_11_en & ram_1_MPORT_11_mask) begin
      ram_1[ram_1_MPORT_11_addr] <= ram_1_MPORT_11_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_12_en & ram_1_MPORT_12_mask) begin
      ram_1[ram_1_MPORT_12_addr] <= ram_1_MPORT_12_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_13_en & ram_1_MPORT_13_mask) begin
      ram_1[ram_1_MPORT_13_addr] <= ram_1_MPORT_13_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_14_en & ram_1_MPORT_14_mask) begin
      ram_1[ram_1_MPORT_14_addr] <= ram_1_MPORT_14_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_15_en & ram_1_MPORT_15_mask) begin
      ram_1[ram_1_MPORT_15_addr] <= ram_1_MPORT_15_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_16_en & ram_1_MPORT_16_mask) begin
      ram_1[ram_1_MPORT_16_addr] <= ram_1_MPORT_16_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_17_en & ram_1_MPORT_17_mask) begin
      ram_1[ram_1_MPORT_17_addr] <= ram_1_MPORT_17_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_18_en & ram_1_MPORT_18_mask) begin
      ram_1[ram_1_MPORT_18_addr] <= ram_1_MPORT_18_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_19_en & ram_1_MPORT_19_mask) begin
      ram_1[ram_1_MPORT_19_addr] <= ram_1_MPORT_19_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_20_en & ram_1_MPORT_20_mask) begin
      ram_1[ram_1_MPORT_20_addr] <= ram_1_MPORT_20_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_21_en & ram_1_MPORT_21_mask) begin
      ram_1[ram_1_MPORT_21_addr] <= ram_1_MPORT_21_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_22_en & ram_1_MPORT_22_mask) begin
      ram_1[ram_1_MPORT_22_addr] <= ram_1_MPORT_22_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_23_en & ram_1_MPORT_23_mask) begin
      ram_1[ram_1_MPORT_23_addr] <= ram_1_MPORT_23_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_24_en & ram_1_MPORT_24_mask) begin
      ram_1[ram_1_MPORT_24_addr] <= ram_1_MPORT_24_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_25_en & ram_1_MPORT_25_mask) begin
      ram_1[ram_1_MPORT_25_addr] <= ram_1_MPORT_25_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_26_en & ram_1_MPORT_26_mask) begin
      ram_1[ram_1_MPORT_26_addr] <= ram_1_MPORT_26_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_27_en & ram_1_MPORT_27_mask) begin
      ram_1[ram_1_MPORT_27_addr] <= ram_1_MPORT_27_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_28_en & ram_1_MPORT_28_mask) begin
      ram_1[ram_1_MPORT_28_addr] <= ram_1_MPORT_28_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_29_en & ram_1_MPORT_29_mask) begin
      ram_1[ram_1_MPORT_29_addr] <= ram_1_MPORT_29_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_30_en & ram_1_MPORT_30_mask) begin
      ram_1[ram_1_MPORT_30_addr] <= ram_1_MPORT_30_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_31_en & ram_1_MPORT_31_mask) begin
      ram_1[ram_1_MPORT_31_addr] <= ram_1_MPORT_31_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_32_en & ram_1_MPORT_32_mask) begin
      ram_1[ram_1_MPORT_32_addr] <= ram_1_MPORT_32_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_33_en & ram_1_MPORT_33_mask) begin
      ram_1[ram_1_MPORT_33_addr] <= ram_1_MPORT_33_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_34_en & ram_1_MPORT_34_mask) begin
      ram_1[ram_1_MPORT_34_addr] <= ram_1_MPORT_34_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_35_en & ram_1_MPORT_35_mask) begin
      ram_1[ram_1_MPORT_35_addr] <= ram_1_MPORT_35_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_36_en & ram_1_MPORT_36_mask) begin
      ram_1[ram_1_MPORT_36_addr] <= ram_1_MPORT_36_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_37_en & ram_1_MPORT_37_mask) begin
      ram_1[ram_1_MPORT_37_addr] <= ram_1_MPORT_37_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_38_en & ram_1_MPORT_38_mask) begin
      ram_1[ram_1_MPORT_38_addr] <= ram_1_MPORT_38_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_39_en & ram_1_MPORT_39_mask) begin
      ram_1[ram_1_MPORT_39_addr] <= ram_1_MPORT_39_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_40_en & ram_1_MPORT_40_mask) begin
      ram_1[ram_1_MPORT_40_addr] <= ram_1_MPORT_40_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_41_en & ram_1_MPORT_41_mask) begin
      ram_1[ram_1_MPORT_41_addr] <= ram_1_MPORT_41_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_42_en & ram_1_MPORT_42_mask) begin
      ram_1[ram_1_MPORT_42_addr] <= ram_1_MPORT_42_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_43_en & ram_1_MPORT_43_mask) begin
      ram_1[ram_1_MPORT_43_addr] <= ram_1_MPORT_43_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_44_en & ram_1_MPORT_44_mask) begin
      ram_1[ram_1_MPORT_44_addr] <= ram_1_MPORT_44_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_45_en & ram_1_MPORT_45_mask) begin
      ram_1[ram_1_MPORT_45_addr] <= ram_1_MPORT_45_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_46_en & ram_1_MPORT_46_mask) begin
      ram_1[ram_1_MPORT_46_addr] <= ram_1_MPORT_46_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_47_en & ram_1_MPORT_47_mask) begin
      ram_1[ram_1_MPORT_47_addr] <= ram_1_MPORT_47_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_48_en & ram_1_MPORT_48_mask) begin
      ram_1[ram_1_MPORT_48_addr] <= ram_1_MPORT_48_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_49_en & ram_1_MPORT_49_mask) begin
      ram_1[ram_1_MPORT_49_addr] <= ram_1_MPORT_49_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_50_en & ram_1_MPORT_50_mask) begin
      ram_1[ram_1_MPORT_50_addr] <= ram_1_MPORT_50_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_51_en & ram_1_MPORT_51_mask) begin
      ram_1[ram_1_MPORT_51_addr] <= ram_1_MPORT_51_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_52_en & ram_1_MPORT_52_mask) begin
      ram_1[ram_1_MPORT_52_addr] <= ram_1_MPORT_52_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_53_en & ram_1_MPORT_53_mask) begin
      ram_1[ram_1_MPORT_53_addr] <= ram_1_MPORT_53_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_54_en & ram_1_MPORT_54_mask) begin
      ram_1[ram_1_MPORT_54_addr] <= ram_1_MPORT_54_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_55_en & ram_1_MPORT_55_mask) begin
      ram_1[ram_1_MPORT_55_addr] <= ram_1_MPORT_55_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_56_en & ram_1_MPORT_56_mask) begin
      ram_1[ram_1_MPORT_56_addr] <= ram_1_MPORT_56_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_57_en & ram_1_MPORT_57_mask) begin
      ram_1[ram_1_MPORT_57_addr] <= ram_1_MPORT_57_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_58_en & ram_1_MPORT_58_mask) begin
      ram_1[ram_1_MPORT_58_addr] <= ram_1_MPORT_58_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_59_en & ram_1_MPORT_59_mask) begin
      ram_1[ram_1_MPORT_59_addr] <= ram_1_MPORT_59_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_60_en & ram_1_MPORT_60_mask) begin
      ram_1[ram_1_MPORT_60_addr] <= ram_1_MPORT_60_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_61_en & ram_1_MPORT_61_mask) begin
      ram_1[ram_1_MPORT_61_addr] <= ram_1_MPORT_61_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_62_en & ram_1_MPORT_62_mask) begin
      ram_1[ram_1_MPORT_62_addr] <= ram_1_MPORT_62_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_63_en & ram_1_MPORT_63_mask) begin
      ram_1[ram_1_MPORT_63_addr] <= ram_1_MPORT_63_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_64_en & ram_1_MPORT_64_mask) begin
      ram_1[ram_1_MPORT_64_addr] <= ram_1_MPORT_64_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_65_en & ram_1_MPORT_65_mask) begin
      ram_1[ram_1_MPORT_65_addr] <= ram_1_MPORT_65_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_66_en & ram_1_MPORT_66_mask) begin
      ram_1[ram_1_MPORT_66_addr] <= ram_1_MPORT_66_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_67_en & ram_1_MPORT_67_mask) begin
      ram_1[ram_1_MPORT_67_addr] <= ram_1_MPORT_67_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_68_en & ram_1_MPORT_68_mask) begin
      ram_1[ram_1_MPORT_68_addr] <= ram_1_MPORT_68_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_69_en & ram_1_MPORT_69_mask) begin
      ram_1[ram_1_MPORT_69_addr] <= ram_1_MPORT_69_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_70_en & ram_1_MPORT_70_mask) begin
      ram_1[ram_1_MPORT_70_addr] <= ram_1_MPORT_70_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_71_en & ram_1_MPORT_71_mask) begin
      ram_1[ram_1_MPORT_71_addr] <= ram_1_MPORT_71_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_72_en & ram_1_MPORT_72_mask) begin
      ram_1[ram_1_MPORT_72_addr] <= ram_1_MPORT_72_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_73_en & ram_1_MPORT_73_mask) begin
      ram_1[ram_1_MPORT_73_addr] <= ram_1_MPORT_73_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_74_en & ram_1_MPORT_74_mask) begin
      ram_1[ram_1_MPORT_74_addr] <= ram_1_MPORT_74_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_75_en & ram_1_MPORT_75_mask) begin
      ram_1[ram_1_MPORT_75_addr] <= ram_1_MPORT_75_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_76_en & ram_1_MPORT_76_mask) begin
      ram_1[ram_1_MPORT_76_addr] <= ram_1_MPORT_76_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_77_en & ram_1_MPORT_77_mask) begin
      ram_1[ram_1_MPORT_77_addr] <= ram_1_MPORT_77_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_78_en & ram_1_MPORT_78_mask) begin
      ram_1[ram_1_MPORT_78_addr] <= ram_1_MPORT_78_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_79_en & ram_1_MPORT_79_mask) begin
      ram_1[ram_1_MPORT_79_addr] <= ram_1_MPORT_79_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_80_en & ram_1_MPORT_80_mask) begin
      ram_1[ram_1_MPORT_80_addr] <= ram_1_MPORT_80_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_81_en & ram_1_MPORT_81_mask) begin
      ram_1[ram_1_MPORT_81_addr] <= ram_1_MPORT_81_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_82_en & ram_1_MPORT_82_mask) begin
      ram_1[ram_1_MPORT_82_addr] <= ram_1_MPORT_82_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_83_en & ram_1_MPORT_83_mask) begin
      ram_1[ram_1_MPORT_83_addr] <= ram_1_MPORT_83_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_84_en & ram_1_MPORT_84_mask) begin
      ram_1[ram_1_MPORT_84_addr] <= ram_1_MPORT_84_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_85_en & ram_1_MPORT_85_mask) begin
      ram_1[ram_1_MPORT_85_addr] <= ram_1_MPORT_85_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_86_en & ram_1_MPORT_86_mask) begin
      ram_1[ram_1_MPORT_86_addr] <= ram_1_MPORT_86_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_87_en & ram_1_MPORT_87_mask) begin
      ram_1[ram_1_MPORT_87_addr] <= ram_1_MPORT_87_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_88_en & ram_1_MPORT_88_mask) begin
      ram_1[ram_1_MPORT_88_addr] <= ram_1_MPORT_88_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_89_en & ram_1_MPORT_89_mask) begin
      ram_1[ram_1_MPORT_89_addr] <= ram_1_MPORT_89_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_90_en & ram_1_MPORT_90_mask) begin
      ram_1[ram_1_MPORT_90_addr] <= ram_1_MPORT_90_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_91_en & ram_1_MPORT_91_mask) begin
      ram_1[ram_1_MPORT_91_addr] <= ram_1_MPORT_91_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_92_en & ram_1_MPORT_92_mask) begin
      ram_1[ram_1_MPORT_92_addr] <= ram_1_MPORT_92_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_93_en & ram_1_MPORT_93_mask) begin
      ram_1[ram_1_MPORT_93_addr] <= ram_1_MPORT_93_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_94_en & ram_1_MPORT_94_mask) begin
      ram_1[ram_1_MPORT_94_addr] <= ram_1_MPORT_94_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_95_en & ram_1_MPORT_95_mask) begin
      ram_1[ram_1_MPORT_95_addr] <= ram_1_MPORT_95_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_96_en & ram_1_MPORT_96_mask) begin
      ram_1[ram_1_MPORT_96_addr] <= ram_1_MPORT_96_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_97_en & ram_1_MPORT_97_mask) begin
      ram_1[ram_1_MPORT_97_addr] <= ram_1_MPORT_97_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_98_en & ram_1_MPORT_98_mask) begin
      ram_1[ram_1_MPORT_98_addr] <= ram_1_MPORT_98_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_99_en & ram_1_MPORT_99_mask) begin
      ram_1[ram_1_MPORT_99_addr] <= ram_1_MPORT_99_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_100_en & ram_1_MPORT_100_mask) begin
      ram_1[ram_1_MPORT_100_addr] <= ram_1_MPORT_100_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_101_en & ram_1_MPORT_101_mask) begin
      ram_1[ram_1_MPORT_101_addr] <= ram_1_MPORT_101_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_102_en & ram_1_MPORT_102_mask) begin
      ram_1[ram_1_MPORT_102_addr] <= ram_1_MPORT_102_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_103_en & ram_1_MPORT_103_mask) begin
      ram_1[ram_1_MPORT_103_addr] <= ram_1_MPORT_103_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_104_en & ram_1_MPORT_104_mask) begin
      ram_1[ram_1_MPORT_104_addr] <= ram_1_MPORT_104_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_105_en & ram_1_MPORT_105_mask) begin
      ram_1[ram_1_MPORT_105_addr] <= ram_1_MPORT_105_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_106_en & ram_1_MPORT_106_mask) begin
      ram_1[ram_1_MPORT_106_addr] <= ram_1_MPORT_106_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_107_en & ram_1_MPORT_107_mask) begin
      ram_1[ram_1_MPORT_107_addr] <= ram_1_MPORT_107_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_108_en & ram_1_MPORT_108_mask) begin
      ram_1[ram_1_MPORT_108_addr] <= ram_1_MPORT_108_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_109_en & ram_1_MPORT_109_mask) begin
      ram_1[ram_1_MPORT_109_addr] <= ram_1_MPORT_109_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_110_en & ram_1_MPORT_110_mask) begin
      ram_1[ram_1_MPORT_110_addr] <= ram_1_MPORT_110_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_111_en & ram_1_MPORT_111_mask) begin
      ram_1[ram_1_MPORT_111_addr] <= ram_1_MPORT_111_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_112_en & ram_1_MPORT_112_mask) begin
      ram_1[ram_1_MPORT_112_addr] <= ram_1_MPORT_112_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_113_en & ram_1_MPORT_113_mask) begin
      ram_1[ram_1_MPORT_113_addr] <= ram_1_MPORT_113_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_114_en & ram_1_MPORT_114_mask) begin
      ram_1[ram_1_MPORT_114_addr] <= ram_1_MPORT_114_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_115_en & ram_1_MPORT_115_mask) begin
      ram_1[ram_1_MPORT_115_addr] <= ram_1_MPORT_115_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_116_en & ram_1_MPORT_116_mask) begin
      ram_1[ram_1_MPORT_116_addr] <= ram_1_MPORT_116_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_117_en & ram_1_MPORT_117_mask) begin
      ram_1[ram_1_MPORT_117_addr] <= ram_1_MPORT_117_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_118_en & ram_1_MPORT_118_mask) begin
      ram_1[ram_1_MPORT_118_addr] <= ram_1_MPORT_118_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_119_en & ram_1_MPORT_119_mask) begin
      ram_1[ram_1_MPORT_119_addr] <= ram_1_MPORT_119_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_120_en & ram_1_MPORT_120_mask) begin
      ram_1[ram_1_MPORT_120_addr] <= ram_1_MPORT_120_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_121_en & ram_1_MPORT_121_mask) begin
      ram_1[ram_1_MPORT_121_addr] <= ram_1_MPORT_121_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_122_en & ram_1_MPORT_122_mask) begin
      ram_1[ram_1_MPORT_122_addr] <= ram_1_MPORT_122_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_123_en & ram_1_MPORT_123_mask) begin
      ram_1[ram_1_MPORT_123_addr] <= ram_1_MPORT_123_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_124_en & ram_1_MPORT_124_mask) begin
      ram_1[ram_1_MPORT_124_addr] <= ram_1_MPORT_124_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_125_en & ram_1_MPORT_125_mask) begin
      ram_1[ram_1_MPORT_125_addr] <= ram_1_MPORT_125_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_126_en & ram_1_MPORT_126_mask) begin
      ram_1[ram_1_MPORT_126_addr] <= ram_1_MPORT_126_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_127_en & ram_1_MPORT_127_mask) begin
      ram_1[ram_1_MPORT_127_addr] <= ram_1_MPORT_127_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_128_en & ram_1_MPORT_128_mask) begin
      ram_1[ram_1_MPORT_128_addr] <= ram_1_MPORT_128_data; // @[SRAM.scala 36:26]
    end
    if (io_rw) begin
      ram_1_io_rdata_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      ram_1_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    end
    if (io_rw ? 1'h0 : 1'h1) begin
      ram_1_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
    if (ram_2_MPORT_en & ram_2_MPORT_mask) begin
      ram_2[ram_2_MPORT_addr] <= ram_2_MPORT_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_1_en & ram_2_MPORT_1_mask) begin
      ram_2[ram_2_MPORT_1_addr] <= ram_2_MPORT_1_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_2_en & ram_2_MPORT_2_mask) begin
      ram_2[ram_2_MPORT_2_addr] <= ram_2_MPORT_2_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_3_en & ram_2_MPORT_3_mask) begin
      ram_2[ram_2_MPORT_3_addr] <= ram_2_MPORT_3_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_4_en & ram_2_MPORT_4_mask) begin
      ram_2[ram_2_MPORT_4_addr] <= ram_2_MPORT_4_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_5_en & ram_2_MPORT_5_mask) begin
      ram_2[ram_2_MPORT_5_addr] <= ram_2_MPORT_5_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_6_en & ram_2_MPORT_6_mask) begin
      ram_2[ram_2_MPORT_6_addr] <= ram_2_MPORT_6_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_7_en & ram_2_MPORT_7_mask) begin
      ram_2[ram_2_MPORT_7_addr] <= ram_2_MPORT_7_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_8_en & ram_2_MPORT_8_mask) begin
      ram_2[ram_2_MPORT_8_addr] <= ram_2_MPORT_8_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_9_en & ram_2_MPORT_9_mask) begin
      ram_2[ram_2_MPORT_9_addr] <= ram_2_MPORT_9_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_10_en & ram_2_MPORT_10_mask) begin
      ram_2[ram_2_MPORT_10_addr] <= ram_2_MPORT_10_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_11_en & ram_2_MPORT_11_mask) begin
      ram_2[ram_2_MPORT_11_addr] <= ram_2_MPORT_11_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_12_en & ram_2_MPORT_12_mask) begin
      ram_2[ram_2_MPORT_12_addr] <= ram_2_MPORT_12_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_13_en & ram_2_MPORT_13_mask) begin
      ram_2[ram_2_MPORT_13_addr] <= ram_2_MPORT_13_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_14_en & ram_2_MPORT_14_mask) begin
      ram_2[ram_2_MPORT_14_addr] <= ram_2_MPORT_14_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_15_en & ram_2_MPORT_15_mask) begin
      ram_2[ram_2_MPORT_15_addr] <= ram_2_MPORT_15_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_16_en & ram_2_MPORT_16_mask) begin
      ram_2[ram_2_MPORT_16_addr] <= ram_2_MPORT_16_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_17_en & ram_2_MPORT_17_mask) begin
      ram_2[ram_2_MPORT_17_addr] <= ram_2_MPORT_17_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_18_en & ram_2_MPORT_18_mask) begin
      ram_2[ram_2_MPORT_18_addr] <= ram_2_MPORT_18_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_19_en & ram_2_MPORT_19_mask) begin
      ram_2[ram_2_MPORT_19_addr] <= ram_2_MPORT_19_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_20_en & ram_2_MPORT_20_mask) begin
      ram_2[ram_2_MPORT_20_addr] <= ram_2_MPORT_20_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_21_en & ram_2_MPORT_21_mask) begin
      ram_2[ram_2_MPORT_21_addr] <= ram_2_MPORT_21_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_22_en & ram_2_MPORT_22_mask) begin
      ram_2[ram_2_MPORT_22_addr] <= ram_2_MPORT_22_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_23_en & ram_2_MPORT_23_mask) begin
      ram_2[ram_2_MPORT_23_addr] <= ram_2_MPORT_23_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_24_en & ram_2_MPORT_24_mask) begin
      ram_2[ram_2_MPORT_24_addr] <= ram_2_MPORT_24_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_25_en & ram_2_MPORT_25_mask) begin
      ram_2[ram_2_MPORT_25_addr] <= ram_2_MPORT_25_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_26_en & ram_2_MPORT_26_mask) begin
      ram_2[ram_2_MPORT_26_addr] <= ram_2_MPORT_26_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_27_en & ram_2_MPORT_27_mask) begin
      ram_2[ram_2_MPORT_27_addr] <= ram_2_MPORT_27_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_28_en & ram_2_MPORT_28_mask) begin
      ram_2[ram_2_MPORT_28_addr] <= ram_2_MPORT_28_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_29_en & ram_2_MPORT_29_mask) begin
      ram_2[ram_2_MPORT_29_addr] <= ram_2_MPORT_29_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_30_en & ram_2_MPORT_30_mask) begin
      ram_2[ram_2_MPORT_30_addr] <= ram_2_MPORT_30_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_31_en & ram_2_MPORT_31_mask) begin
      ram_2[ram_2_MPORT_31_addr] <= ram_2_MPORT_31_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_32_en & ram_2_MPORT_32_mask) begin
      ram_2[ram_2_MPORT_32_addr] <= ram_2_MPORT_32_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_33_en & ram_2_MPORT_33_mask) begin
      ram_2[ram_2_MPORT_33_addr] <= ram_2_MPORT_33_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_34_en & ram_2_MPORT_34_mask) begin
      ram_2[ram_2_MPORT_34_addr] <= ram_2_MPORT_34_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_35_en & ram_2_MPORT_35_mask) begin
      ram_2[ram_2_MPORT_35_addr] <= ram_2_MPORT_35_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_36_en & ram_2_MPORT_36_mask) begin
      ram_2[ram_2_MPORT_36_addr] <= ram_2_MPORT_36_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_37_en & ram_2_MPORT_37_mask) begin
      ram_2[ram_2_MPORT_37_addr] <= ram_2_MPORT_37_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_38_en & ram_2_MPORT_38_mask) begin
      ram_2[ram_2_MPORT_38_addr] <= ram_2_MPORT_38_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_39_en & ram_2_MPORT_39_mask) begin
      ram_2[ram_2_MPORT_39_addr] <= ram_2_MPORT_39_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_40_en & ram_2_MPORT_40_mask) begin
      ram_2[ram_2_MPORT_40_addr] <= ram_2_MPORT_40_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_41_en & ram_2_MPORT_41_mask) begin
      ram_2[ram_2_MPORT_41_addr] <= ram_2_MPORT_41_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_42_en & ram_2_MPORT_42_mask) begin
      ram_2[ram_2_MPORT_42_addr] <= ram_2_MPORT_42_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_43_en & ram_2_MPORT_43_mask) begin
      ram_2[ram_2_MPORT_43_addr] <= ram_2_MPORT_43_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_44_en & ram_2_MPORT_44_mask) begin
      ram_2[ram_2_MPORT_44_addr] <= ram_2_MPORT_44_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_45_en & ram_2_MPORT_45_mask) begin
      ram_2[ram_2_MPORT_45_addr] <= ram_2_MPORT_45_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_46_en & ram_2_MPORT_46_mask) begin
      ram_2[ram_2_MPORT_46_addr] <= ram_2_MPORT_46_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_47_en & ram_2_MPORT_47_mask) begin
      ram_2[ram_2_MPORT_47_addr] <= ram_2_MPORT_47_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_48_en & ram_2_MPORT_48_mask) begin
      ram_2[ram_2_MPORT_48_addr] <= ram_2_MPORT_48_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_49_en & ram_2_MPORT_49_mask) begin
      ram_2[ram_2_MPORT_49_addr] <= ram_2_MPORT_49_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_50_en & ram_2_MPORT_50_mask) begin
      ram_2[ram_2_MPORT_50_addr] <= ram_2_MPORT_50_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_51_en & ram_2_MPORT_51_mask) begin
      ram_2[ram_2_MPORT_51_addr] <= ram_2_MPORT_51_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_52_en & ram_2_MPORT_52_mask) begin
      ram_2[ram_2_MPORT_52_addr] <= ram_2_MPORT_52_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_53_en & ram_2_MPORT_53_mask) begin
      ram_2[ram_2_MPORT_53_addr] <= ram_2_MPORT_53_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_54_en & ram_2_MPORT_54_mask) begin
      ram_2[ram_2_MPORT_54_addr] <= ram_2_MPORT_54_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_55_en & ram_2_MPORT_55_mask) begin
      ram_2[ram_2_MPORT_55_addr] <= ram_2_MPORT_55_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_56_en & ram_2_MPORT_56_mask) begin
      ram_2[ram_2_MPORT_56_addr] <= ram_2_MPORT_56_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_57_en & ram_2_MPORT_57_mask) begin
      ram_2[ram_2_MPORT_57_addr] <= ram_2_MPORT_57_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_58_en & ram_2_MPORT_58_mask) begin
      ram_2[ram_2_MPORT_58_addr] <= ram_2_MPORT_58_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_59_en & ram_2_MPORT_59_mask) begin
      ram_2[ram_2_MPORT_59_addr] <= ram_2_MPORT_59_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_60_en & ram_2_MPORT_60_mask) begin
      ram_2[ram_2_MPORT_60_addr] <= ram_2_MPORT_60_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_61_en & ram_2_MPORT_61_mask) begin
      ram_2[ram_2_MPORT_61_addr] <= ram_2_MPORT_61_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_62_en & ram_2_MPORT_62_mask) begin
      ram_2[ram_2_MPORT_62_addr] <= ram_2_MPORT_62_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_63_en & ram_2_MPORT_63_mask) begin
      ram_2[ram_2_MPORT_63_addr] <= ram_2_MPORT_63_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_64_en & ram_2_MPORT_64_mask) begin
      ram_2[ram_2_MPORT_64_addr] <= ram_2_MPORT_64_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_65_en & ram_2_MPORT_65_mask) begin
      ram_2[ram_2_MPORT_65_addr] <= ram_2_MPORT_65_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_66_en & ram_2_MPORT_66_mask) begin
      ram_2[ram_2_MPORT_66_addr] <= ram_2_MPORT_66_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_67_en & ram_2_MPORT_67_mask) begin
      ram_2[ram_2_MPORT_67_addr] <= ram_2_MPORT_67_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_68_en & ram_2_MPORT_68_mask) begin
      ram_2[ram_2_MPORT_68_addr] <= ram_2_MPORT_68_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_69_en & ram_2_MPORT_69_mask) begin
      ram_2[ram_2_MPORT_69_addr] <= ram_2_MPORT_69_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_70_en & ram_2_MPORT_70_mask) begin
      ram_2[ram_2_MPORT_70_addr] <= ram_2_MPORT_70_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_71_en & ram_2_MPORT_71_mask) begin
      ram_2[ram_2_MPORT_71_addr] <= ram_2_MPORT_71_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_72_en & ram_2_MPORT_72_mask) begin
      ram_2[ram_2_MPORT_72_addr] <= ram_2_MPORT_72_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_73_en & ram_2_MPORT_73_mask) begin
      ram_2[ram_2_MPORT_73_addr] <= ram_2_MPORT_73_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_74_en & ram_2_MPORT_74_mask) begin
      ram_2[ram_2_MPORT_74_addr] <= ram_2_MPORT_74_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_75_en & ram_2_MPORT_75_mask) begin
      ram_2[ram_2_MPORT_75_addr] <= ram_2_MPORT_75_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_76_en & ram_2_MPORT_76_mask) begin
      ram_2[ram_2_MPORT_76_addr] <= ram_2_MPORT_76_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_77_en & ram_2_MPORT_77_mask) begin
      ram_2[ram_2_MPORT_77_addr] <= ram_2_MPORT_77_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_78_en & ram_2_MPORT_78_mask) begin
      ram_2[ram_2_MPORT_78_addr] <= ram_2_MPORT_78_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_79_en & ram_2_MPORT_79_mask) begin
      ram_2[ram_2_MPORT_79_addr] <= ram_2_MPORT_79_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_80_en & ram_2_MPORT_80_mask) begin
      ram_2[ram_2_MPORT_80_addr] <= ram_2_MPORT_80_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_81_en & ram_2_MPORT_81_mask) begin
      ram_2[ram_2_MPORT_81_addr] <= ram_2_MPORT_81_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_82_en & ram_2_MPORT_82_mask) begin
      ram_2[ram_2_MPORT_82_addr] <= ram_2_MPORT_82_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_83_en & ram_2_MPORT_83_mask) begin
      ram_2[ram_2_MPORT_83_addr] <= ram_2_MPORT_83_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_84_en & ram_2_MPORT_84_mask) begin
      ram_2[ram_2_MPORT_84_addr] <= ram_2_MPORT_84_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_85_en & ram_2_MPORT_85_mask) begin
      ram_2[ram_2_MPORT_85_addr] <= ram_2_MPORT_85_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_86_en & ram_2_MPORT_86_mask) begin
      ram_2[ram_2_MPORT_86_addr] <= ram_2_MPORT_86_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_87_en & ram_2_MPORT_87_mask) begin
      ram_2[ram_2_MPORT_87_addr] <= ram_2_MPORT_87_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_88_en & ram_2_MPORT_88_mask) begin
      ram_2[ram_2_MPORT_88_addr] <= ram_2_MPORT_88_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_89_en & ram_2_MPORT_89_mask) begin
      ram_2[ram_2_MPORT_89_addr] <= ram_2_MPORT_89_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_90_en & ram_2_MPORT_90_mask) begin
      ram_2[ram_2_MPORT_90_addr] <= ram_2_MPORT_90_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_91_en & ram_2_MPORT_91_mask) begin
      ram_2[ram_2_MPORT_91_addr] <= ram_2_MPORT_91_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_92_en & ram_2_MPORT_92_mask) begin
      ram_2[ram_2_MPORT_92_addr] <= ram_2_MPORT_92_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_93_en & ram_2_MPORT_93_mask) begin
      ram_2[ram_2_MPORT_93_addr] <= ram_2_MPORT_93_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_94_en & ram_2_MPORT_94_mask) begin
      ram_2[ram_2_MPORT_94_addr] <= ram_2_MPORT_94_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_95_en & ram_2_MPORT_95_mask) begin
      ram_2[ram_2_MPORT_95_addr] <= ram_2_MPORT_95_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_96_en & ram_2_MPORT_96_mask) begin
      ram_2[ram_2_MPORT_96_addr] <= ram_2_MPORT_96_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_97_en & ram_2_MPORT_97_mask) begin
      ram_2[ram_2_MPORT_97_addr] <= ram_2_MPORT_97_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_98_en & ram_2_MPORT_98_mask) begin
      ram_2[ram_2_MPORT_98_addr] <= ram_2_MPORT_98_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_99_en & ram_2_MPORT_99_mask) begin
      ram_2[ram_2_MPORT_99_addr] <= ram_2_MPORT_99_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_100_en & ram_2_MPORT_100_mask) begin
      ram_2[ram_2_MPORT_100_addr] <= ram_2_MPORT_100_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_101_en & ram_2_MPORT_101_mask) begin
      ram_2[ram_2_MPORT_101_addr] <= ram_2_MPORT_101_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_102_en & ram_2_MPORT_102_mask) begin
      ram_2[ram_2_MPORT_102_addr] <= ram_2_MPORT_102_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_103_en & ram_2_MPORT_103_mask) begin
      ram_2[ram_2_MPORT_103_addr] <= ram_2_MPORT_103_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_104_en & ram_2_MPORT_104_mask) begin
      ram_2[ram_2_MPORT_104_addr] <= ram_2_MPORT_104_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_105_en & ram_2_MPORT_105_mask) begin
      ram_2[ram_2_MPORT_105_addr] <= ram_2_MPORT_105_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_106_en & ram_2_MPORT_106_mask) begin
      ram_2[ram_2_MPORT_106_addr] <= ram_2_MPORT_106_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_107_en & ram_2_MPORT_107_mask) begin
      ram_2[ram_2_MPORT_107_addr] <= ram_2_MPORT_107_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_108_en & ram_2_MPORT_108_mask) begin
      ram_2[ram_2_MPORT_108_addr] <= ram_2_MPORT_108_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_109_en & ram_2_MPORT_109_mask) begin
      ram_2[ram_2_MPORT_109_addr] <= ram_2_MPORT_109_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_110_en & ram_2_MPORT_110_mask) begin
      ram_2[ram_2_MPORT_110_addr] <= ram_2_MPORT_110_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_111_en & ram_2_MPORT_111_mask) begin
      ram_2[ram_2_MPORT_111_addr] <= ram_2_MPORT_111_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_112_en & ram_2_MPORT_112_mask) begin
      ram_2[ram_2_MPORT_112_addr] <= ram_2_MPORT_112_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_113_en & ram_2_MPORT_113_mask) begin
      ram_2[ram_2_MPORT_113_addr] <= ram_2_MPORT_113_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_114_en & ram_2_MPORT_114_mask) begin
      ram_2[ram_2_MPORT_114_addr] <= ram_2_MPORT_114_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_115_en & ram_2_MPORT_115_mask) begin
      ram_2[ram_2_MPORT_115_addr] <= ram_2_MPORT_115_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_116_en & ram_2_MPORT_116_mask) begin
      ram_2[ram_2_MPORT_116_addr] <= ram_2_MPORT_116_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_117_en & ram_2_MPORT_117_mask) begin
      ram_2[ram_2_MPORT_117_addr] <= ram_2_MPORT_117_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_118_en & ram_2_MPORT_118_mask) begin
      ram_2[ram_2_MPORT_118_addr] <= ram_2_MPORT_118_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_119_en & ram_2_MPORT_119_mask) begin
      ram_2[ram_2_MPORT_119_addr] <= ram_2_MPORT_119_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_120_en & ram_2_MPORT_120_mask) begin
      ram_2[ram_2_MPORT_120_addr] <= ram_2_MPORT_120_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_121_en & ram_2_MPORT_121_mask) begin
      ram_2[ram_2_MPORT_121_addr] <= ram_2_MPORT_121_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_122_en & ram_2_MPORT_122_mask) begin
      ram_2[ram_2_MPORT_122_addr] <= ram_2_MPORT_122_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_123_en & ram_2_MPORT_123_mask) begin
      ram_2[ram_2_MPORT_123_addr] <= ram_2_MPORT_123_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_124_en & ram_2_MPORT_124_mask) begin
      ram_2[ram_2_MPORT_124_addr] <= ram_2_MPORT_124_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_125_en & ram_2_MPORT_125_mask) begin
      ram_2[ram_2_MPORT_125_addr] <= ram_2_MPORT_125_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_126_en & ram_2_MPORT_126_mask) begin
      ram_2[ram_2_MPORT_126_addr] <= ram_2_MPORT_126_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_127_en & ram_2_MPORT_127_mask) begin
      ram_2[ram_2_MPORT_127_addr] <= ram_2_MPORT_127_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_128_en & ram_2_MPORT_128_mask) begin
      ram_2[ram_2_MPORT_128_addr] <= ram_2_MPORT_128_data; // @[SRAM.scala 36:26]
    end
    if (io_rw) begin
      ram_2_io_rdata_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      ram_2_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    end
    if (io_rw ? 1'h0 : 1'h1) begin
      ram_2_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
    if (ram_3_MPORT_en & ram_3_MPORT_mask) begin
      ram_3[ram_3_MPORT_addr] <= ram_3_MPORT_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_1_en & ram_3_MPORT_1_mask) begin
      ram_3[ram_3_MPORT_1_addr] <= ram_3_MPORT_1_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_2_en & ram_3_MPORT_2_mask) begin
      ram_3[ram_3_MPORT_2_addr] <= ram_3_MPORT_2_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_3_en & ram_3_MPORT_3_mask) begin
      ram_3[ram_3_MPORT_3_addr] <= ram_3_MPORT_3_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_4_en & ram_3_MPORT_4_mask) begin
      ram_3[ram_3_MPORT_4_addr] <= ram_3_MPORT_4_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_5_en & ram_3_MPORT_5_mask) begin
      ram_3[ram_3_MPORT_5_addr] <= ram_3_MPORT_5_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_6_en & ram_3_MPORT_6_mask) begin
      ram_3[ram_3_MPORT_6_addr] <= ram_3_MPORT_6_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_7_en & ram_3_MPORT_7_mask) begin
      ram_3[ram_3_MPORT_7_addr] <= ram_3_MPORT_7_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_8_en & ram_3_MPORT_8_mask) begin
      ram_3[ram_3_MPORT_8_addr] <= ram_3_MPORT_8_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_9_en & ram_3_MPORT_9_mask) begin
      ram_3[ram_3_MPORT_9_addr] <= ram_3_MPORT_9_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_10_en & ram_3_MPORT_10_mask) begin
      ram_3[ram_3_MPORT_10_addr] <= ram_3_MPORT_10_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_11_en & ram_3_MPORT_11_mask) begin
      ram_3[ram_3_MPORT_11_addr] <= ram_3_MPORT_11_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_12_en & ram_3_MPORT_12_mask) begin
      ram_3[ram_3_MPORT_12_addr] <= ram_3_MPORT_12_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_13_en & ram_3_MPORT_13_mask) begin
      ram_3[ram_3_MPORT_13_addr] <= ram_3_MPORT_13_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_14_en & ram_3_MPORT_14_mask) begin
      ram_3[ram_3_MPORT_14_addr] <= ram_3_MPORT_14_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_15_en & ram_3_MPORT_15_mask) begin
      ram_3[ram_3_MPORT_15_addr] <= ram_3_MPORT_15_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_16_en & ram_3_MPORT_16_mask) begin
      ram_3[ram_3_MPORT_16_addr] <= ram_3_MPORT_16_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_17_en & ram_3_MPORT_17_mask) begin
      ram_3[ram_3_MPORT_17_addr] <= ram_3_MPORT_17_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_18_en & ram_3_MPORT_18_mask) begin
      ram_3[ram_3_MPORT_18_addr] <= ram_3_MPORT_18_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_19_en & ram_3_MPORT_19_mask) begin
      ram_3[ram_3_MPORT_19_addr] <= ram_3_MPORT_19_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_20_en & ram_3_MPORT_20_mask) begin
      ram_3[ram_3_MPORT_20_addr] <= ram_3_MPORT_20_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_21_en & ram_3_MPORT_21_mask) begin
      ram_3[ram_3_MPORT_21_addr] <= ram_3_MPORT_21_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_22_en & ram_3_MPORT_22_mask) begin
      ram_3[ram_3_MPORT_22_addr] <= ram_3_MPORT_22_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_23_en & ram_3_MPORT_23_mask) begin
      ram_3[ram_3_MPORT_23_addr] <= ram_3_MPORT_23_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_24_en & ram_3_MPORT_24_mask) begin
      ram_3[ram_3_MPORT_24_addr] <= ram_3_MPORT_24_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_25_en & ram_3_MPORT_25_mask) begin
      ram_3[ram_3_MPORT_25_addr] <= ram_3_MPORT_25_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_26_en & ram_3_MPORT_26_mask) begin
      ram_3[ram_3_MPORT_26_addr] <= ram_3_MPORT_26_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_27_en & ram_3_MPORT_27_mask) begin
      ram_3[ram_3_MPORT_27_addr] <= ram_3_MPORT_27_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_28_en & ram_3_MPORT_28_mask) begin
      ram_3[ram_3_MPORT_28_addr] <= ram_3_MPORT_28_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_29_en & ram_3_MPORT_29_mask) begin
      ram_3[ram_3_MPORT_29_addr] <= ram_3_MPORT_29_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_30_en & ram_3_MPORT_30_mask) begin
      ram_3[ram_3_MPORT_30_addr] <= ram_3_MPORT_30_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_31_en & ram_3_MPORT_31_mask) begin
      ram_3[ram_3_MPORT_31_addr] <= ram_3_MPORT_31_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_32_en & ram_3_MPORT_32_mask) begin
      ram_3[ram_3_MPORT_32_addr] <= ram_3_MPORT_32_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_33_en & ram_3_MPORT_33_mask) begin
      ram_3[ram_3_MPORT_33_addr] <= ram_3_MPORT_33_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_34_en & ram_3_MPORT_34_mask) begin
      ram_3[ram_3_MPORT_34_addr] <= ram_3_MPORT_34_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_35_en & ram_3_MPORT_35_mask) begin
      ram_3[ram_3_MPORT_35_addr] <= ram_3_MPORT_35_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_36_en & ram_3_MPORT_36_mask) begin
      ram_3[ram_3_MPORT_36_addr] <= ram_3_MPORT_36_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_37_en & ram_3_MPORT_37_mask) begin
      ram_3[ram_3_MPORT_37_addr] <= ram_3_MPORT_37_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_38_en & ram_3_MPORT_38_mask) begin
      ram_3[ram_3_MPORT_38_addr] <= ram_3_MPORT_38_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_39_en & ram_3_MPORT_39_mask) begin
      ram_3[ram_3_MPORT_39_addr] <= ram_3_MPORT_39_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_40_en & ram_3_MPORT_40_mask) begin
      ram_3[ram_3_MPORT_40_addr] <= ram_3_MPORT_40_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_41_en & ram_3_MPORT_41_mask) begin
      ram_3[ram_3_MPORT_41_addr] <= ram_3_MPORT_41_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_42_en & ram_3_MPORT_42_mask) begin
      ram_3[ram_3_MPORT_42_addr] <= ram_3_MPORT_42_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_43_en & ram_3_MPORT_43_mask) begin
      ram_3[ram_3_MPORT_43_addr] <= ram_3_MPORT_43_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_44_en & ram_3_MPORT_44_mask) begin
      ram_3[ram_3_MPORT_44_addr] <= ram_3_MPORT_44_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_45_en & ram_3_MPORT_45_mask) begin
      ram_3[ram_3_MPORT_45_addr] <= ram_3_MPORT_45_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_46_en & ram_3_MPORT_46_mask) begin
      ram_3[ram_3_MPORT_46_addr] <= ram_3_MPORT_46_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_47_en & ram_3_MPORT_47_mask) begin
      ram_3[ram_3_MPORT_47_addr] <= ram_3_MPORT_47_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_48_en & ram_3_MPORT_48_mask) begin
      ram_3[ram_3_MPORT_48_addr] <= ram_3_MPORT_48_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_49_en & ram_3_MPORT_49_mask) begin
      ram_3[ram_3_MPORT_49_addr] <= ram_3_MPORT_49_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_50_en & ram_3_MPORT_50_mask) begin
      ram_3[ram_3_MPORT_50_addr] <= ram_3_MPORT_50_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_51_en & ram_3_MPORT_51_mask) begin
      ram_3[ram_3_MPORT_51_addr] <= ram_3_MPORT_51_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_52_en & ram_3_MPORT_52_mask) begin
      ram_3[ram_3_MPORT_52_addr] <= ram_3_MPORT_52_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_53_en & ram_3_MPORT_53_mask) begin
      ram_3[ram_3_MPORT_53_addr] <= ram_3_MPORT_53_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_54_en & ram_3_MPORT_54_mask) begin
      ram_3[ram_3_MPORT_54_addr] <= ram_3_MPORT_54_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_55_en & ram_3_MPORT_55_mask) begin
      ram_3[ram_3_MPORT_55_addr] <= ram_3_MPORT_55_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_56_en & ram_3_MPORT_56_mask) begin
      ram_3[ram_3_MPORT_56_addr] <= ram_3_MPORT_56_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_57_en & ram_3_MPORT_57_mask) begin
      ram_3[ram_3_MPORT_57_addr] <= ram_3_MPORT_57_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_58_en & ram_3_MPORT_58_mask) begin
      ram_3[ram_3_MPORT_58_addr] <= ram_3_MPORT_58_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_59_en & ram_3_MPORT_59_mask) begin
      ram_3[ram_3_MPORT_59_addr] <= ram_3_MPORT_59_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_60_en & ram_3_MPORT_60_mask) begin
      ram_3[ram_3_MPORT_60_addr] <= ram_3_MPORT_60_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_61_en & ram_3_MPORT_61_mask) begin
      ram_3[ram_3_MPORT_61_addr] <= ram_3_MPORT_61_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_62_en & ram_3_MPORT_62_mask) begin
      ram_3[ram_3_MPORT_62_addr] <= ram_3_MPORT_62_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_63_en & ram_3_MPORT_63_mask) begin
      ram_3[ram_3_MPORT_63_addr] <= ram_3_MPORT_63_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_64_en & ram_3_MPORT_64_mask) begin
      ram_3[ram_3_MPORT_64_addr] <= ram_3_MPORT_64_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_65_en & ram_3_MPORT_65_mask) begin
      ram_3[ram_3_MPORT_65_addr] <= ram_3_MPORT_65_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_66_en & ram_3_MPORT_66_mask) begin
      ram_3[ram_3_MPORT_66_addr] <= ram_3_MPORT_66_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_67_en & ram_3_MPORT_67_mask) begin
      ram_3[ram_3_MPORT_67_addr] <= ram_3_MPORT_67_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_68_en & ram_3_MPORT_68_mask) begin
      ram_3[ram_3_MPORT_68_addr] <= ram_3_MPORT_68_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_69_en & ram_3_MPORT_69_mask) begin
      ram_3[ram_3_MPORT_69_addr] <= ram_3_MPORT_69_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_70_en & ram_3_MPORT_70_mask) begin
      ram_3[ram_3_MPORT_70_addr] <= ram_3_MPORT_70_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_71_en & ram_3_MPORT_71_mask) begin
      ram_3[ram_3_MPORT_71_addr] <= ram_3_MPORT_71_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_72_en & ram_3_MPORT_72_mask) begin
      ram_3[ram_3_MPORT_72_addr] <= ram_3_MPORT_72_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_73_en & ram_3_MPORT_73_mask) begin
      ram_3[ram_3_MPORT_73_addr] <= ram_3_MPORT_73_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_74_en & ram_3_MPORT_74_mask) begin
      ram_3[ram_3_MPORT_74_addr] <= ram_3_MPORT_74_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_75_en & ram_3_MPORT_75_mask) begin
      ram_3[ram_3_MPORT_75_addr] <= ram_3_MPORT_75_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_76_en & ram_3_MPORT_76_mask) begin
      ram_3[ram_3_MPORT_76_addr] <= ram_3_MPORT_76_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_77_en & ram_3_MPORT_77_mask) begin
      ram_3[ram_3_MPORT_77_addr] <= ram_3_MPORT_77_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_78_en & ram_3_MPORT_78_mask) begin
      ram_3[ram_3_MPORT_78_addr] <= ram_3_MPORT_78_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_79_en & ram_3_MPORT_79_mask) begin
      ram_3[ram_3_MPORT_79_addr] <= ram_3_MPORT_79_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_80_en & ram_3_MPORT_80_mask) begin
      ram_3[ram_3_MPORT_80_addr] <= ram_3_MPORT_80_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_81_en & ram_3_MPORT_81_mask) begin
      ram_3[ram_3_MPORT_81_addr] <= ram_3_MPORT_81_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_82_en & ram_3_MPORT_82_mask) begin
      ram_3[ram_3_MPORT_82_addr] <= ram_3_MPORT_82_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_83_en & ram_3_MPORT_83_mask) begin
      ram_3[ram_3_MPORT_83_addr] <= ram_3_MPORT_83_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_84_en & ram_3_MPORT_84_mask) begin
      ram_3[ram_3_MPORT_84_addr] <= ram_3_MPORT_84_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_85_en & ram_3_MPORT_85_mask) begin
      ram_3[ram_3_MPORT_85_addr] <= ram_3_MPORT_85_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_86_en & ram_3_MPORT_86_mask) begin
      ram_3[ram_3_MPORT_86_addr] <= ram_3_MPORT_86_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_87_en & ram_3_MPORT_87_mask) begin
      ram_3[ram_3_MPORT_87_addr] <= ram_3_MPORT_87_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_88_en & ram_3_MPORT_88_mask) begin
      ram_3[ram_3_MPORT_88_addr] <= ram_3_MPORT_88_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_89_en & ram_3_MPORT_89_mask) begin
      ram_3[ram_3_MPORT_89_addr] <= ram_3_MPORT_89_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_90_en & ram_3_MPORT_90_mask) begin
      ram_3[ram_3_MPORT_90_addr] <= ram_3_MPORT_90_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_91_en & ram_3_MPORT_91_mask) begin
      ram_3[ram_3_MPORT_91_addr] <= ram_3_MPORT_91_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_92_en & ram_3_MPORT_92_mask) begin
      ram_3[ram_3_MPORT_92_addr] <= ram_3_MPORT_92_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_93_en & ram_3_MPORT_93_mask) begin
      ram_3[ram_3_MPORT_93_addr] <= ram_3_MPORT_93_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_94_en & ram_3_MPORT_94_mask) begin
      ram_3[ram_3_MPORT_94_addr] <= ram_3_MPORT_94_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_95_en & ram_3_MPORT_95_mask) begin
      ram_3[ram_3_MPORT_95_addr] <= ram_3_MPORT_95_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_96_en & ram_3_MPORT_96_mask) begin
      ram_3[ram_3_MPORT_96_addr] <= ram_3_MPORT_96_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_97_en & ram_3_MPORT_97_mask) begin
      ram_3[ram_3_MPORT_97_addr] <= ram_3_MPORT_97_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_98_en & ram_3_MPORT_98_mask) begin
      ram_3[ram_3_MPORT_98_addr] <= ram_3_MPORT_98_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_99_en & ram_3_MPORT_99_mask) begin
      ram_3[ram_3_MPORT_99_addr] <= ram_3_MPORT_99_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_100_en & ram_3_MPORT_100_mask) begin
      ram_3[ram_3_MPORT_100_addr] <= ram_3_MPORT_100_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_101_en & ram_3_MPORT_101_mask) begin
      ram_3[ram_3_MPORT_101_addr] <= ram_3_MPORT_101_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_102_en & ram_3_MPORT_102_mask) begin
      ram_3[ram_3_MPORT_102_addr] <= ram_3_MPORT_102_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_103_en & ram_3_MPORT_103_mask) begin
      ram_3[ram_3_MPORT_103_addr] <= ram_3_MPORT_103_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_104_en & ram_3_MPORT_104_mask) begin
      ram_3[ram_3_MPORT_104_addr] <= ram_3_MPORT_104_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_105_en & ram_3_MPORT_105_mask) begin
      ram_3[ram_3_MPORT_105_addr] <= ram_3_MPORT_105_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_106_en & ram_3_MPORT_106_mask) begin
      ram_3[ram_3_MPORT_106_addr] <= ram_3_MPORT_106_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_107_en & ram_3_MPORT_107_mask) begin
      ram_3[ram_3_MPORT_107_addr] <= ram_3_MPORT_107_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_108_en & ram_3_MPORT_108_mask) begin
      ram_3[ram_3_MPORT_108_addr] <= ram_3_MPORT_108_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_109_en & ram_3_MPORT_109_mask) begin
      ram_3[ram_3_MPORT_109_addr] <= ram_3_MPORT_109_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_110_en & ram_3_MPORT_110_mask) begin
      ram_3[ram_3_MPORT_110_addr] <= ram_3_MPORT_110_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_111_en & ram_3_MPORT_111_mask) begin
      ram_3[ram_3_MPORT_111_addr] <= ram_3_MPORT_111_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_112_en & ram_3_MPORT_112_mask) begin
      ram_3[ram_3_MPORT_112_addr] <= ram_3_MPORT_112_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_113_en & ram_3_MPORT_113_mask) begin
      ram_3[ram_3_MPORT_113_addr] <= ram_3_MPORT_113_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_114_en & ram_3_MPORT_114_mask) begin
      ram_3[ram_3_MPORT_114_addr] <= ram_3_MPORT_114_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_115_en & ram_3_MPORT_115_mask) begin
      ram_3[ram_3_MPORT_115_addr] <= ram_3_MPORT_115_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_116_en & ram_3_MPORT_116_mask) begin
      ram_3[ram_3_MPORT_116_addr] <= ram_3_MPORT_116_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_117_en & ram_3_MPORT_117_mask) begin
      ram_3[ram_3_MPORT_117_addr] <= ram_3_MPORT_117_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_118_en & ram_3_MPORT_118_mask) begin
      ram_3[ram_3_MPORT_118_addr] <= ram_3_MPORT_118_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_119_en & ram_3_MPORT_119_mask) begin
      ram_3[ram_3_MPORT_119_addr] <= ram_3_MPORT_119_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_120_en & ram_3_MPORT_120_mask) begin
      ram_3[ram_3_MPORT_120_addr] <= ram_3_MPORT_120_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_121_en & ram_3_MPORT_121_mask) begin
      ram_3[ram_3_MPORT_121_addr] <= ram_3_MPORT_121_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_122_en & ram_3_MPORT_122_mask) begin
      ram_3[ram_3_MPORT_122_addr] <= ram_3_MPORT_122_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_123_en & ram_3_MPORT_123_mask) begin
      ram_3[ram_3_MPORT_123_addr] <= ram_3_MPORT_123_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_124_en & ram_3_MPORT_124_mask) begin
      ram_3[ram_3_MPORT_124_addr] <= ram_3_MPORT_124_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_125_en & ram_3_MPORT_125_mask) begin
      ram_3[ram_3_MPORT_125_addr] <= ram_3_MPORT_125_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_126_en & ram_3_MPORT_126_mask) begin
      ram_3[ram_3_MPORT_126_addr] <= ram_3_MPORT_126_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_127_en & ram_3_MPORT_127_mask) begin
      ram_3[ram_3_MPORT_127_addr] <= ram_3_MPORT_127_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_128_en & ram_3_MPORT_128_mask) begin
      ram_3[ram_3_MPORT_128_addr] <= ram_3_MPORT_128_data; // @[SRAM.scala 36:26]
    end
    if (io_rw) begin
      ram_3_io_rdata_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      ram_3_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    end
    if (io_rw ? 1'h0 : 1'h1) begin
      ram_3_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_0[initvar] = _RAND_0[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_1[initvar] = _RAND_3[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_2[initvar] = _RAND_6[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_3[initvar] = _RAND_9[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_0_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_0_io_rdata_MPORT_addr_pipe_0 = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  ram_1_io_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ram_1_io_rdata_MPORT_addr_pipe_0 = _RAND_5[6:0];
  _RAND_7 = {1{`RANDOM}};
  ram_2_io_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ram_2_io_rdata_MPORT_addr_pipe_0 = _RAND_8[6:0];
  _RAND_10 = {1{`RANDOM}};
  ram_3_io_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ram_3_io_rdata_MPORT_addr_pipe_0 = _RAND_11[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
