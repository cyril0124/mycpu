module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_inst,
  input         io_enq_bits_valid,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_inst,
  output        io_deq_bits_valid,
  output [3:0]  io_count,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_inst [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_inst_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_inst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_inst_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_inst_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_inst_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_inst_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_inst_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_valid [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_valid_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_valid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_valid_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_valid_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_valid_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_valid_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_valid_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [2:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 326:32]
  wire [3:0] _io_count_T_1 = maybe_full & ptr_match ? 4'h8 : 4'h0; // @[Decoupled.scala 329:20]
  wire [3:0] _GEN_12 = {{1'd0}, ptr_diff}; // @[Decoupled.scala 329:62]
  assign ram_inst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_inst_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_inst_io_deq_bits_MPORT_data = ram_inst[ram_inst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_inst_MPORT_data = io_enq_bits_inst;
  assign ram_inst_MPORT_addr = enq_ptr_value;
  assign ram_inst_MPORT_mask = 1'h1;
  assign ram_inst_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_valid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_valid_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_valid_io_deq_bits_MPORT_data = ram_valid[ram_valid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_valid_MPORT_data = io_enq_bits_valid;
  assign ram_valid_MPORT_addr = enq_ptr_value;
  assign ram_valid_MPORT_mask = 1'h1;
  assign ram_valid_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_inst = ram_inst_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_valid = ram_valid_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_count = _io_count_T_1 | _GEN_12; // @[Decoupled.scala 329:62]
  always @(posedge clock) begin
    if (ram_inst_MPORT_en & ram_inst_MPORT_mask) begin
      ram_inst[ram_inst_MPORT_addr] <= ram_inst_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_valid_MPORT_en & ram_valid_MPORT_mask) begin
      ram_valid[ram_valid_MPORT_addr] <= ram_valid_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      enq_ptr_value <= 3'h0; // @[Counter.scala 98:11]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      deq_ptr_value <= 3'h0; // @[Counter.scala 98:11]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      maybe_full <= 1'h0; // @[Decoupled.scala 299:16]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_inst[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_valid[initvar] = _RAND_1[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      enq_ptr_value <= 3'h0; // @[Counter.scala 98:11]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      deq_ptr_value <= 3'h0; // @[Counter.scala 98:11]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      maybe_full <= 1'h0; // @[Decoupled.scala 299:16]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstBuffer(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_icache_data,
  input  [31:0] io_in_bits_icache_addr,
  input  [31:0] io_in_bits_icache_inst_0,
  input  [31:0] io_in_bits_icache_inst_1,
  input  [31:0] io_in_bits_icache_inst_2,
  input  [31:0] io_in_bits_icache_inst_3,
  input  [2:0]  io_in_bits_icache_size,
  input  [31:0] io_in_bits_pc,
  input         io_in_bits_flush,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_inst_0_inst,
  output        io_out_bits_inst_0_valid,
  output [31:0] io_out_bits_inst_1_inst,
  output        io_out_bits_inst_1_valid,
  output [31:0] io_out_bits_inst_2_inst,
  output        io_out_bits_inst_2_valid,
  output [31:0] io_out_bits_inst_3_inst,
  output        io_out_bits_inst_3_valid,
  output [31:0] io_out_bits_pc,
  output        io_status_back_pressure,
  output        io_status_full
);
  wire  entries_0_clock; // @[InstBuffer.scala 37:48]
  wire  entries_0_reset; // @[InstBuffer.scala 37:48]
  wire  entries_0_io_enq_ready; // @[InstBuffer.scala 37:48]
  wire  entries_0_io_enq_valid; // @[InstBuffer.scala 37:48]
  wire [31:0] entries_0_io_enq_bits_inst; // @[InstBuffer.scala 37:48]
  wire  entries_0_io_enq_bits_valid; // @[InstBuffer.scala 37:48]
  wire  entries_0_io_deq_ready; // @[InstBuffer.scala 37:48]
  wire  entries_0_io_deq_valid; // @[InstBuffer.scala 37:48]
  wire [31:0] entries_0_io_deq_bits_inst; // @[InstBuffer.scala 37:48]
  wire  entries_0_io_deq_bits_valid; // @[InstBuffer.scala 37:48]
  wire [3:0] entries_0_io_count; // @[InstBuffer.scala 37:48]
  wire  entries_0_io_flush; // @[InstBuffer.scala 37:48]
  wire  entries_1_clock; // @[InstBuffer.scala 37:48]
  wire  entries_1_reset; // @[InstBuffer.scala 37:48]
  wire  entries_1_io_enq_ready; // @[InstBuffer.scala 37:48]
  wire  entries_1_io_enq_valid; // @[InstBuffer.scala 37:48]
  wire [31:0] entries_1_io_enq_bits_inst; // @[InstBuffer.scala 37:48]
  wire  entries_1_io_enq_bits_valid; // @[InstBuffer.scala 37:48]
  wire  entries_1_io_deq_ready; // @[InstBuffer.scala 37:48]
  wire  entries_1_io_deq_valid; // @[InstBuffer.scala 37:48]
  wire [31:0] entries_1_io_deq_bits_inst; // @[InstBuffer.scala 37:48]
  wire  entries_1_io_deq_bits_valid; // @[InstBuffer.scala 37:48]
  wire [3:0] entries_1_io_count; // @[InstBuffer.scala 37:48]
  wire  entries_1_io_flush; // @[InstBuffer.scala 37:48]
  wire  entries_2_clock; // @[InstBuffer.scala 37:48]
  wire  entries_2_reset; // @[InstBuffer.scala 37:48]
  wire  entries_2_io_enq_ready; // @[InstBuffer.scala 37:48]
  wire  entries_2_io_enq_valid; // @[InstBuffer.scala 37:48]
  wire [31:0] entries_2_io_enq_bits_inst; // @[InstBuffer.scala 37:48]
  wire  entries_2_io_enq_bits_valid; // @[InstBuffer.scala 37:48]
  wire  entries_2_io_deq_ready; // @[InstBuffer.scala 37:48]
  wire  entries_2_io_deq_valid; // @[InstBuffer.scala 37:48]
  wire [31:0] entries_2_io_deq_bits_inst; // @[InstBuffer.scala 37:48]
  wire  entries_2_io_deq_bits_valid; // @[InstBuffer.scala 37:48]
  wire [3:0] entries_2_io_count; // @[InstBuffer.scala 37:48]
  wire  entries_2_io_flush; // @[InstBuffer.scala 37:48]
  wire  entries_3_clock; // @[InstBuffer.scala 37:48]
  wire  entries_3_reset; // @[InstBuffer.scala 37:48]
  wire  entries_3_io_enq_ready; // @[InstBuffer.scala 37:48]
  wire  entries_3_io_enq_valid; // @[InstBuffer.scala 37:48]
  wire [31:0] entries_3_io_enq_bits_inst; // @[InstBuffer.scala 37:48]
  wire  entries_3_io_enq_bits_valid; // @[InstBuffer.scala 37:48]
  wire  entries_3_io_deq_ready; // @[InstBuffer.scala 37:48]
  wire  entries_3_io_deq_valid; // @[InstBuffer.scala 37:48]
  wire [31:0] entries_3_io_deq_bits_inst; // @[InstBuffer.scala 37:48]
  wire  entries_3_io_deq_bits_valid; // @[InstBuffer.scala 37:48]
  wire [3:0] entries_3_io_count; // @[InstBuffer.scala 37:48]
  wire  entries_3_io_flush; // @[InstBuffer.scala 37:48]
  wire  pcQueue_clock; // @[InstBuffer.scala 38:25]
  wire  pcQueue_reset; // @[InstBuffer.scala 38:25]
  wire  pcQueue_io_enq_ready; // @[InstBuffer.scala 38:25]
  wire  pcQueue_io_enq_valid; // @[InstBuffer.scala 38:25]
  wire [31:0] pcQueue_io_enq_bits; // @[InstBuffer.scala 38:25]
  wire  pcQueue_io_deq_ready; // @[InstBuffer.scala 38:25]
  wire  pcQueue_io_deq_valid; // @[InstBuffer.scala 38:25]
  wire [31:0] pcQueue_io_deq_bits; // @[InstBuffer.scala 38:25]
  wire  pcQueue_io_flush; // @[InstBuffer.scala 38:25]
  wire [2:0] _mask_T_2 = 3'h4 - io_in_bits_icache_size; // @[InstBuffer.scala 46:56]
  wire [3:0] mask = 4'hf >> _mask_T_2; // @[InstBuffer.scala 46:37]
  Queue entries_0 ( // @[InstBuffer.scala 37:48]
    .clock(entries_0_clock),
    .reset(entries_0_reset),
    .io_enq_ready(entries_0_io_enq_ready),
    .io_enq_valid(entries_0_io_enq_valid),
    .io_enq_bits_inst(entries_0_io_enq_bits_inst),
    .io_enq_bits_valid(entries_0_io_enq_bits_valid),
    .io_deq_ready(entries_0_io_deq_ready),
    .io_deq_valid(entries_0_io_deq_valid),
    .io_deq_bits_inst(entries_0_io_deq_bits_inst),
    .io_deq_bits_valid(entries_0_io_deq_bits_valid),
    .io_count(entries_0_io_count),
    .io_flush(entries_0_io_flush)
  );
  Queue entries_1 ( // @[InstBuffer.scala 37:48]
    .clock(entries_1_clock),
    .reset(entries_1_reset),
    .io_enq_ready(entries_1_io_enq_ready),
    .io_enq_valid(entries_1_io_enq_valid),
    .io_enq_bits_inst(entries_1_io_enq_bits_inst),
    .io_enq_bits_valid(entries_1_io_enq_bits_valid),
    .io_deq_ready(entries_1_io_deq_ready),
    .io_deq_valid(entries_1_io_deq_valid),
    .io_deq_bits_inst(entries_1_io_deq_bits_inst),
    .io_deq_bits_valid(entries_1_io_deq_bits_valid),
    .io_count(entries_1_io_count),
    .io_flush(entries_1_io_flush)
  );
  Queue entries_2 ( // @[InstBuffer.scala 37:48]
    .clock(entries_2_clock),
    .reset(entries_2_reset),
    .io_enq_ready(entries_2_io_enq_ready),
    .io_enq_valid(entries_2_io_enq_valid),
    .io_enq_bits_inst(entries_2_io_enq_bits_inst),
    .io_enq_bits_valid(entries_2_io_enq_bits_valid),
    .io_deq_ready(entries_2_io_deq_ready),
    .io_deq_valid(entries_2_io_deq_valid),
    .io_deq_bits_inst(entries_2_io_deq_bits_inst),
    .io_deq_bits_valid(entries_2_io_deq_bits_valid),
    .io_count(entries_2_io_count),
    .io_flush(entries_2_io_flush)
  );
  Queue entries_3 ( // @[InstBuffer.scala 37:48]
    .clock(entries_3_clock),
    .reset(entries_3_reset),
    .io_enq_ready(entries_3_io_enq_ready),
    .io_enq_valid(entries_3_io_enq_valid),
    .io_enq_bits_inst(entries_3_io_enq_bits_inst),
    .io_enq_bits_valid(entries_3_io_enq_bits_valid),
    .io_deq_ready(entries_3_io_deq_ready),
    .io_deq_valid(entries_3_io_deq_valid),
    .io_deq_bits_inst(entries_3_io_deq_bits_inst),
    .io_deq_bits_valid(entries_3_io_deq_bits_valid),
    .io_count(entries_3_io_count),
    .io_flush(entries_3_io_flush)
  );
  Queue_4 pcQueue ( // @[InstBuffer.scala 38:25]
    .clock(pcQueue_clock),
    .reset(pcQueue_reset),
    .io_enq_ready(pcQueue_io_enq_ready),
    .io_enq_valid(pcQueue_io_enq_valid),
    .io_enq_bits(pcQueue_io_enq_bits),
    .io_deq_ready(pcQueue_io_deq_ready),
    .io_deq_valid(pcQueue_io_deq_valid),
    .io_deq_bits(pcQueue_io_deq_bits),
    .io_flush(pcQueue_io_flush)
  );
  assign io_in_ready = entries_0_io_enq_ready & entries_1_io_enq_ready & entries_2_io_enq_ready & entries_3_io_enq_ready
    ; // @[InstBuffer.scala 42:61]
  assign io_out_valid = entries_0_io_deq_valid & entries_1_io_deq_valid & entries_2_io_deq_valid &
    entries_3_io_deq_valid; // @[InstBuffer.scala 43:62]
  assign io_out_bits_inst_0_inst = entries_0_io_deq_bits_inst; // @[InstBuffer.scala 53:29]
  assign io_out_bits_inst_0_valid = entries_0_io_deq_bits_valid; // @[InstBuffer.scala 53:29]
  assign io_out_bits_inst_1_inst = entries_1_io_deq_bits_inst; // @[InstBuffer.scala 53:29]
  assign io_out_bits_inst_1_valid = entries_1_io_deq_bits_valid; // @[InstBuffer.scala 53:29]
  assign io_out_bits_inst_2_inst = entries_2_io_deq_bits_inst; // @[InstBuffer.scala 53:29]
  assign io_out_bits_inst_2_valid = entries_2_io_deq_bits_valid; // @[InstBuffer.scala 53:29]
  assign io_out_bits_inst_3_inst = entries_3_io_deq_bits_inst; // @[InstBuffer.scala 53:29]
  assign io_out_bits_inst_3_valid = entries_3_io_deq_bits_valid; // @[InstBuffer.scala 53:29]
  assign io_out_bits_pc = pcQueue_io_deq_bits; // @[InstBuffer.scala 60:20]
  assign io_status_back_pressure = entries_0_io_count >= 4'h5; // @[InstBuffer.scala 40:52]
  assign io_status_full = entries_0_io_count == 4'h6; // @[InstBuffer.scala 41:43]
  assign entries_0_clock = clock;
  assign entries_0_reset = reset;
  assign entries_0_io_enq_valid = io_in_valid; // @[InstBuffer.scala 49:33]
  assign entries_0_io_enq_bits_inst = io_in_bits_icache_inst_0; // @[InstBuffer.scala 50:37]
  assign entries_0_io_enq_bits_valid = mask[0]; // @[InstBuffer.scala 51:45]
  assign entries_0_io_deq_ready = io_out_ready; // @[InstBuffer.scala 52:33]
  assign entries_0_io_flush = io_in_bits_flush; // @[InstBuffer.scala 48:33]
  assign entries_1_clock = clock;
  assign entries_1_reset = reset;
  assign entries_1_io_enq_valid = io_in_valid; // @[InstBuffer.scala 49:33]
  assign entries_1_io_enq_bits_inst = io_in_bits_icache_inst_1; // @[InstBuffer.scala 50:37]
  assign entries_1_io_enq_bits_valid = mask[1]; // @[InstBuffer.scala 51:45]
  assign entries_1_io_deq_ready = io_out_ready; // @[InstBuffer.scala 52:33]
  assign entries_1_io_flush = io_in_bits_flush; // @[InstBuffer.scala 48:33]
  assign entries_2_clock = clock;
  assign entries_2_reset = reset;
  assign entries_2_io_enq_valid = io_in_valid; // @[InstBuffer.scala 49:33]
  assign entries_2_io_enq_bits_inst = io_in_bits_icache_inst_2; // @[InstBuffer.scala 50:37]
  assign entries_2_io_enq_bits_valid = mask[2]; // @[InstBuffer.scala 51:45]
  assign entries_2_io_deq_ready = io_out_ready; // @[InstBuffer.scala 52:33]
  assign entries_2_io_flush = io_in_bits_flush; // @[InstBuffer.scala 48:33]
  assign entries_3_clock = clock;
  assign entries_3_reset = reset;
  assign entries_3_io_enq_valid = io_in_valid; // @[InstBuffer.scala 49:33]
  assign entries_3_io_enq_bits_inst = io_in_bits_icache_inst_3; // @[InstBuffer.scala 50:37]
  assign entries_3_io_enq_bits_valid = mask[3]; // @[InstBuffer.scala 51:45]
  assign entries_3_io_deq_ready = io_out_ready; // @[InstBuffer.scala 52:33]
  assign entries_3_io_flush = io_in_bits_flush; // @[InstBuffer.scala 48:33]
  assign pcQueue_clock = clock;
  assign pcQueue_reset = reset;
  assign pcQueue_io_enq_valid = io_in_valid; // @[InstBuffer.scala 58:26]
  assign pcQueue_io_enq_bits = io_in_bits_pc; // @[InstBuffer.scala 57:25]
  assign pcQueue_io_deq_ready = io_out_ready; // @[InstBuffer.scala 61:26]
  assign pcQueue_io_flush = io_in_bits_flush; // @[InstBuffer.scala 56:26]
endmodule
module BankRAM_2P(
  input         clock,
  input         reset,
  input  [6:0]  io_r_addr,
  output [31:0] io_r_data,
  input         io_w_en,
  input  [6:0]  io_w_addr,
  input  [31:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:127]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [6:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 32'h0;
  assign mem_MPORT_addr = 7'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 32'h0;
  assign mem_MPORT_1_addr = 7'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 32'h0;
  assign mem_MPORT_2_addr = 7'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 32'h0;
  assign mem_MPORT_3_addr = 7'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 32'h0;
  assign mem_MPORT_4_addr = 7'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 32'h0;
  assign mem_MPORT_5_addr = 7'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 32'h0;
  assign mem_MPORT_6_addr = 7'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 32'h0;
  assign mem_MPORT_7_addr = 7'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 32'h0;
  assign mem_MPORT_8_addr = 7'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 32'h0;
  assign mem_MPORT_9_addr = 7'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 32'h0;
  assign mem_MPORT_10_addr = 7'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 32'h0;
  assign mem_MPORT_11_addr = 7'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 32'h0;
  assign mem_MPORT_12_addr = 7'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 32'h0;
  assign mem_MPORT_13_addr = 7'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 32'h0;
  assign mem_MPORT_14_addr = 7'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 32'h0;
  assign mem_MPORT_15_addr = 7'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 32'h0;
  assign mem_MPORT_16_addr = 7'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 32'h0;
  assign mem_MPORT_17_addr = 7'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 32'h0;
  assign mem_MPORT_18_addr = 7'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 32'h0;
  assign mem_MPORT_19_addr = 7'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 32'h0;
  assign mem_MPORT_20_addr = 7'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 32'h0;
  assign mem_MPORT_21_addr = 7'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 32'h0;
  assign mem_MPORT_22_addr = 7'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 32'h0;
  assign mem_MPORT_23_addr = 7'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 32'h0;
  assign mem_MPORT_24_addr = 7'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 32'h0;
  assign mem_MPORT_25_addr = 7'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 32'h0;
  assign mem_MPORT_26_addr = 7'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 32'h0;
  assign mem_MPORT_27_addr = 7'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 32'h0;
  assign mem_MPORT_28_addr = 7'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 32'h0;
  assign mem_MPORT_29_addr = 7'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 32'h0;
  assign mem_MPORT_30_addr = 7'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 32'h0;
  assign mem_MPORT_31_addr = 7'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 32'h0;
  assign mem_MPORT_32_addr = 7'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 32'h0;
  assign mem_MPORT_33_addr = 7'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 32'h0;
  assign mem_MPORT_34_addr = 7'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 32'h0;
  assign mem_MPORT_35_addr = 7'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 32'h0;
  assign mem_MPORT_36_addr = 7'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 32'h0;
  assign mem_MPORT_37_addr = 7'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 32'h0;
  assign mem_MPORT_38_addr = 7'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 32'h0;
  assign mem_MPORT_39_addr = 7'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 32'h0;
  assign mem_MPORT_40_addr = 7'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 32'h0;
  assign mem_MPORT_41_addr = 7'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 32'h0;
  assign mem_MPORT_42_addr = 7'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 32'h0;
  assign mem_MPORT_43_addr = 7'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 32'h0;
  assign mem_MPORT_44_addr = 7'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 32'h0;
  assign mem_MPORT_45_addr = 7'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 32'h0;
  assign mem_MPORT_46_addr = 7'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 32'h0;
  assign mem_MPORT_47_addr = 7'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 32'h0;
  assign mem_MPORT_48_addr = 7'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 32'h0;
  assign mem_MPORT_49_addr = 7'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 32'h0;
  assign mem_MPORT_50_addr = 7'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 32'h0;
  assign mem_MPORT_51_addr = 7'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 32'h0;
  assign mem_MPORT_52_addr = 7'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 32'h0;
  assign mem_MPORT_53_addr = 7'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 32'h0;
  assign mem_MPORT_54_addr = 7'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 32'h0;
  assign mem_MPORT_55_addr = 7'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 32'h0;
  assign mem_MPORT_56_addr = 7'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 32'h0;
  assign mem_MPORT_57_addr = 7'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 32'h0;
  assign mem_MPORT_58_addr = 7'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 32'h0;
  assign mem_MPORT_59_addr = 7'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 32'h0;
  assign mem_MPORT_60_addr = 7'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 32'h0;
  assign mem_MPORT_61_addr = 7'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 32'h0;
  assign mem_MPORT_62_addr = 7'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 32'h0;
  assign mem_MPORT_63_addr = 7'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 32'h0;
  assign mem_MPORT_64_addr = 7'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 32'h0;
  assign mem_MPORT_65_addr = 7'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 32'h0;
  assign mem_MPORT_66_addr = 7'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 32'h0;
  assign mem_MPORT_67_addr = 7'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 32'h0;
  assign mem_MPORT_68_addr = 7'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 32'h0;
  assign mem_MPORT_69_addr = 7'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 32'h0;
  assign mem_MPORT_70_addr = 7'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 32'h0;
  assign mem_MPORT_71_addr = 7'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 32'h0;
  assign mem_MPORT_72_addr = 7'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 32'h0;
  assign mem_MPORT_73_addr = 7'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 32'h0;
  assign mem_MPORT_74_addr = 7'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 32'h0;
  assign mem_MPORT_75_addr = 7'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 32'h0;
  assign mem_MPORT_76_addr = 7'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 32'h0;
  assign mem_MPORT_77_addr = 7'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 32'h0;
  assign mem_MPORT_78_addr = 7'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 32'h0;
  assign mem_MPORT_79_addr = 7'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 32'h0;
  assign mem_MPORT_80_addr = 7'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 32'h0;
  assign mem_MPORT_81_addr = 7'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 32'h0;
  assign mem_MPORT_82_addr = 7'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 32'h0;
  assign mem_MPORT_83_addr = 7'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 32'h0;
  assign mem_MPORT_84_addr = 7'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 32'h0;
  assign mem_MPORT_85_addr = 7'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 32'h0;
  assign mem_MPORT_86_addr = 7'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 32'h0;
  assign mem_MPORT_87_addr = 7'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 32'h0;
  assign mem_MPORT_88_addr = 7'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 32'h0;
  assign mem_MPORT_89_addr = 7'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 32'h0;
  assign mem_MPORT_90_addr = 7'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 32'h0;
  assign mem_MPORT_91_addr = 7'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 32'h0;
  assign mem_MPORT_92_addr = 7'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 32'h0;
  assign mem_MPORT_93_addr = 7'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 32'h0;
  assign mem_MPORT_94_addr = 7'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 32'h0;
  assign mem_MPORT_95_addr = 7'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 32'h0;
  assign mem_MPORT_96_addr = 7'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 32'h0;
  assign mem_MPORT_97_addr = 7'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 32'h0;
  assign mem_MPORT_98_addr = 7'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 32'h0;
  assign mem_MPORT_99_addr = 7'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 32'h0;
  assign mem_MPORT_100_addr = 7'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 32'h0;
  assign mem_MPORT_101_addr = 7'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 32'h0;
  assign mem_MPORT_102_addr = 7'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 32'h0;
  assign mem_MPORT_103_addr = 7'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 32'h0;
  assign mem_MPORT_104_addr = 7'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 32'h0;
  assign mem_MPORT_105_addr = 7'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 32'h0;
  assign mem_MPORT_106_addr = 7'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 32'h0;
  assign mem_MPORT_107_addr = 7'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 32'h0;
  assign mem_MPORT_108_addr = 7'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 32'h0;
  assign mem_MPORT_109_addr = 7'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 32'h0;
  assign mem_MPORT_110_addr = 7'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 32'h0;
  assign mem_MPORT_111_addr = 7'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 32'h0;
  assign mem_MPORT_112_addr = 7'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 32'h0;
  assign mem_MPORT_113_addr = 7'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 32'h0;
  assign mem_MPORT_114_addr = 7'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 32'h0;
  assign mem_MPORT_115_addr = 7'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 32'h0;
  assign mem_MPORT_116_addr = 7'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 32'h0;
  assign mem_MPORT_117_addr = 7'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 32'h0;
  assign mem_MPORT_118_addr = 7'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 32'h0;
  assign mem_MPORT_119_addr = 7'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 32'h0;
  assign mem_MPORT_120_addr = 7'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 32'h0;
  assign mem_MPORT_121_addr = 7'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 32'h0;
  assign mem_MPORT_122_addr = 7'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 32'h0;
  assign mem_MPORT_123_addr = 7'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 32'h0;
  assign mem_MPORT_124_addr = 7'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 32'h0;
  assign mem_MPORT_125_addr = 7'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 32'h0;
  assign mem_MPORT_126_addr = 7'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 32'h0;
  assign mem_MPORT_127_addr = 7'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = io_w_data;
  assign mem_MPORT_128_addr = io_w_addr;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P(
  input         clock,
  input         reset,
  input  [6:0]  io_r_addr,
  output [31:0] io_r_data_0,
  output [31:0] io_r_data_1,
  output [31:0] io_r_data_2,
  output [31:0] io_r_data_3,
  output [31:0] io_r_data_4,
  output [31:0] io_r_data_5,
  output [31:0] io_r_data_6,
  output [31:0] io_r_data_7,
  input         io_w_en,
  input  [6:0]  io_w_addr,
  input  [31:0] io_w_data_0,
  input  [31:0] io_w_data_1,
  input  [31:0] io_w_data_2,
  input  [31:0] io_w_data_3,
  input  [31:0] io_w_data_4,
  input  [31:0] io_w_data_5,
  input  [31:0] io_w_data_6,
  input  [31:0] io_w_data_7,
  input  [7:0]  io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_clock; // @[SRAM_1.scala 201:38]
  wire  brams_4_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_4_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_4_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_clock; // @[SRAM_1.scala 201:38]
  wire  brams_5_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_5_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_5_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_clock; // @[SRAM_1.scala 201:38]
  wire  brams_6_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_6_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_6_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_clock; // @[SRAM_1.scala 201:38]
  wire  brams_7_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_7_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_7_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  BankRAM_2P brams_4 ( // @[SRAM_1.scala 201:38]
    .clock(brams_4_clock),
    .reset(brams_4_reset),
    .io_r_addr(brams_4_io_r_addr),
    .io_r_data(brams_4_io_r_data),
    .io_w_en(brams_4_io_w_en),
    .io_w_addr(brams_4_io_w_addr),
    .io_w_data(brams_4_io_w_data)
  );
  BankRAM_2P brams_5 ( // @[SRAM_1.scala 201:38]
    .clock(brams_5_clock),
    .reset(brams_5_reset),
    .io_r_addr(brams_5_io_r_addr),
    .io_r_data(brams_5_io_r_data),
    .io_w_en(brams_5_io_w_en),
    .io_w_addr(brams_5_io_w_addr),
    .io_w_data(brams_5_io_w_data)
  );
  BankRAM_2P brams_6 ( // @[SRAM_1.scala 201:38]
    .clock(brams_6_clock),
    .reset(brams_6_reset),
    .io_r_addr(brams_6_io_r_addr),
    .io_r_data(brams_6_io_r_data),
    .io_w_en(brams_6_io_w_en),
    .io_w_addr(brams_6_io_w_addr),
    .io_w_data(brams_6_io_w_data)
  );
  BankRAM_2P brams_7 ( // @[SRAM_1.scala 201:38]
    .clock(brams_7_clock),
    .reset(brams_7_reset),
    .io_r_addr(brams_7_io_r_addr),
    .io_r_data(brams_7_io_r_data),
    .io_w_en(brams_7_io_w_en),
    .io_w_addr(brams_7_io_w_addr),
    .io_w_data(brams_7_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_4 = brams_4_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_5 = brams_5_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_6 = brams_6_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_7 = brams_7_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
  assign brams_4_clock = clock;
  assign brams_4_reset = reset;
  assign brams_4_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_4_io_w_en = io_w_en & io_w_maskOH[4]; // @[SRAM_1.scala 208:37]
  assign brams_4_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_4_io_w_data = io_w_data_4; // @[SRAM_1.scala 210:28]
  assign brams_5_clock = clock;
  assign brams_5_reset = reset;
  assign brams_5_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_5_io_w_en = io_w_en & io_w_maskOH[5]; // @[SRAM_1.scala 208:37]
  assign brams_5_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_5_io_w_data = io_w_data_5; // @[SRAM_1.scala 210:28]
  assign brams_6_clock = clock;
  assign brams_6_reset = reset;
  assign brams_6_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_6_io_w_en = io_w_en & io_w_maskOH[6]; // @[SRAM_1.scala 208:37]
  assign brams_6_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_6_io_w_data = io_w_data_6; // @[SRAM_1.scala 210:28]
  assign brams_7_clock = clock;
  assign brams_7_reset = reset;
  assign brams_7_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_7_io_w_en = io_w_en & io_w_maskOH[7]; // @[SRAM_1.scala 208:37]
  assign brams_7_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_7_io_w_data = io_w_data_7; // @[SRAM_1.scala 210:28]
endmodule
module DataBankArray(
  input         clock,
  input         reset,
  output        io_read_req_ready,
  input         io_read_req_valid,
  input  [6:0]  io_read_req_bits_set,
  output [31:0] io_read_resp_0_0,
  output [31:0] io_read_resp_0_1,
  output [31:0] io_read_resp_0_2,
  output [31:0] io_read_resp_0_3,
  output [31:0] io_read_resp_0_4,
  output [31:0] io_read_resp_0_5,
  output [31:0] io_read_resp_0_6,
  output [31:0] io_read_resp_0_7,
  output [31:0] io_read_resp_1_0,
  output [31:0] io_read_resp_1_1,
  output [31:0] io_read_resp_1_2,
  output [31:0] io_read_resp_1_3,
  output [31:0] io_read_resp_1_4,
  output [31:0] io_read_resp_1_5,
  output [31:0] io_read_resp_1_6,
  output [31:0] io_read_resp_1_7,
  output [31:0] io_read_resp_2_0,
  output [31:0] io_read_resp_2_1,
  output [31:0] io_read_resp_2_2,
  output [31:0] io_read_resp_2_3,
  output [31:0] io_read_resp_2_4,
  output [31:0] io_read_resp_2_5,
  output [31:0] io_read_resp_2_6,
  output [31:0] io_read_resp_2_7,
  output [31:0] io_read_resp_3_0,
  output [31:0] io_read_resp_3_1,
  output [31:0] io_read_resp_3_2,
  output [31:0] io_read_resp_3_3,
  output [31:0] io_read_resp_3_4,
  output [31:0] io_read_resp_3_5,
  output [31:0] io_read_resp_3_6,
  output [31:0] io_read_resp_3_7,
  output [31:0] io_read_resp_4_0,
  output [31:0] io_read_resp_4_1,
  output [31:0] io_read_resp_4_2,
  output [31:0] io_read_resp_4_3,
  output [31:0] io_read_resp_4_4,
  output [31:0] io_read_resp_4_5,
  output [31:0] io_read_resp_4_6,
  output [31:0] io_read_resp_4_7,
  output [31:0] io_read_resp_5_0,
  output [31:0] io_read_resp_5_1,
  output [31:0] io_read_resp_5_2,
  output [31:0] io_read_resp_5_3,
  output [31:0] io_read_resp_5_4,
  output [31:0] io_read_resp_5_5,
  output [31:0] io_read_resp_5_6,
  output [31:0] io_read_resp_5_7,
  output [31:0] io_read_resp_6_0,
  output [31:0] io_read_resp_6_1,
  output [31:0] io_read_resp_6_2,
  output [31:0] io_read_resp_6_3,
  output [31:0] io_read_resp_6_4,
  output [31:0] io_read_resp_6_5,
  output [31:0] io_read_resp_6_6,
  output [31:0] io_read_resp_6_7,
  output [31:0] io_read_resp_7_0,
  output [31:0] io_read_resp_7_1,
  output [31:0] io_read_resp_7_2,
  output [31:0] io_read_resp_7_3,
  output [31:0] io_read_resp_7_4,
  output [31:0] io_read_resp_7_5,
  output [31:0] io_read_resp_7_6,
  output [31:0] io_read_resp_7_7,
  output        io_write_req_ready,
  input         io_write_req_valid,
  input  [6:0]  io_write_req_bits_set,
  input  [31:0] io_write_req_bits_data_0,
  input  [31:0] io_write_req_bits_data_1,
  input  [31:0] io_write_req_bits_data_2,
  input  [31:0] io_write_req_bits_data_3,
  input  [31:0] io_write_req_bits_data_4,
  input  [31:0] io_write_req_bits_data_5,
  input  [31:0] io_write_req_bits_data_6,
  input  [31:0] io_write_req_bits_data_7,
  input  [7:0]  io_write_req_bits_blockMask,
  input  [7:0]  io_write_req_bits_way
);
  wire  dataBanks_0_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_0_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_0_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_0_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_0_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_0_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_1_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_1_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_1_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_2_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_2_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_2_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_3_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_3_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_3_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_4_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_4_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_4_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_4_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_4_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_4_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_5_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_5_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_5_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_5_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_5_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_5_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_6_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_6_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_6_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_6_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_6_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_6_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_7_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_7_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_7_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_7_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_7_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_7_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  ren = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  wire  _wen_T_1 = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  SRAMArray_2P dataBanks_0 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_0_clock),
    .reset(dataBanks_0_reset),
    .io_r_addr(dataBanks_0_io_r_addr),
    .io_r_data_0(dataBanks_0_io_r_data_0),
    .io_r_data_1(dataBanks_0_io_r_data_1),
    .io_r_data_2(dataBanks_0_io_r_data_2),
    .io_r_data_3(dataBanks_0_io_r_data_3),
    .io_r_data_4(dataBanks_0_io_r_data_4),
    .io_r_data_5(dataBanks_0_io_r_data_5),
    .io_r_data_6(dataBanks_0_io_r_data_6),
    .io_r_data_7(dataBanks_0_io_r_data_7),
    .io_w_en(dataBanks_0_io_w_en),
    .io_w_addr(dataBanks_0_io_w_addr),
    .io_w_data_0(dataBanks_0_io_w_data_0),
    .io_w_data_1(dataBanks_0_io_w_data_1),
    .io_w_data_2(dataBanks_0_io_w_data_2),
    .io_w_data_3(dataBanks_0_io_w_data_3),
    .io_w_data_4(dataBanks_0_io_w_data_4),
    .io_w_data_5(dataBanks_0_io_w_data_5),
    .io_w_data_6(dataBanks_0_io_w_data_6),
    .io_w_data_7(dataBanks_0_io_w_data_7),
    .io_w_maskOH(dataBanks_0_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_1 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_1_clock),
    .reset(dataBanks_1_reset),
    .io_r_addr(dataBanks_1_io_r_addr),
    .io_r_data_0(dataBanks_1_io_r_data_0),
    .io_r_data_1(dataBanks_1_io_r_data_1),
    .io_r_data_2(dataBanks_1_io_r_data_2),
    .io_r_data_3(dataBanks_1_io_r_data_3),
    .io_r_data_4(dataBanks_1_io_r_data_4),
    .io_r_data_5(dataBanks_1_io_r_data_5),
    .io_r_data_6(dataBanks_1_io_r_data_6),
    .io_r_data_7(dataBanks_1_io_r_data_7),
    .io_w_en(dataBanks_1_io_w_en),
    .io_w_addr(dataBanks_1_io_w_addr),
    .io_w_data_0(dataBanks_1_io_w_data_0),
    .io_w_data_1(dataBanks_1_io_w_data_1),
    .io_w_data_2(dataBanks_1_io_w_data_2),
    .io_w_data_3(dataBanks_1_io_w_data_3),
    .io_w_data_4(dataBanks_1_io_w_data_4),
    .io_w_data_5(dataBanks_1_io_w_data_5),
    .io_w_data_6(dataBanks_1_io_w_data_6),
    .io_w_data_7(dataBanks_1_io_w_data_7),
    .io_w_maskOH(dataBanks_1_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_2 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_2_clock),
    .reset(dataBanks_2_reset),
    .io_r_addr(dataBanks_2_io_r_addr),
    .io_r_data_0(dataBanks_2_io_r_data_0),
    .io_r_data_1(dataBanks_2_io_r_data_1),
    .io_r_data_2(dataBanks_2_io_r_data_2),
    .io_r_data_3(dataBanks_2_io_r_data_3),
    .io_r_data_4(dataBanks_2_io_r_data_4),
    .io_r_data_5(dataBanks_2_io_r_data_5),
    .io_r_data_6(dataBanks_2_io_r_data_6),
    .io_r_data_7(dataBanks_2_io_r_data_7),
    .io_w_en(dataBanks_2_io_w_en),
    .io_w_addr(dataBanks_2_io_w_addr),
    .io_w_data_0(dataBanks_2_io_w_data_0),
    .io_w_data_1(dataBanks_2_io_w_data_1),
    .io_w_data_2(dataBanks_2_io_w_data_2),
    .io_w_data_3(dataBanks_2_io_w_data_3),
    .io_w_data_4(dataBanks_2_io_w_data_4),
    .io_w_data_5(dataBanks_2_io_w_data_5),
    .io_w_data_6(dataBanks_2_io_w_data_6),
    .io_w_data_7(dataBanks_2_io_w_data_7),
    .io_w_maskOH(dataBanks_2_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_3 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_3_clock),
    .reset(dataBanks_3_reset),
    .io_r_addr(dataBanks_3_io_r_addr),
    .io_r_data_0(dataBanks_3_io_r_data_0),
    .io_r_data_1(dataBanks_3_io_r_data_1),
    .io_r_data_2(dataBanks_3_io_r_data_2),
    .io_r_data_3(dataBanks_3_io_r_data_3),
    .io_r_data_4(dataBanks_3_io_r_data_4),
    .io_r_data_5(dataBanks_3_io_r_data_5),
    .io_r_data_6(dataBanks_3_io_r_data_6),
    .io_r_data_7(dataBanks_3_io_r_data_7),
    .io_w_en(dataBanks_3_io_w_en),
    .io_w_addr(dataBanks_3_io_w_addr),
    .io_w_data_0(dataBanks_3_io_w_data_0),
    .io_w_data_1(dataBanks_3_io_w_data_1),
    .io_w_data_2(dataBanks_3_io_w_data_2),
    .io_w_data_3(dataBanks_3_io_w_data_3),
    .io_w_data_4(dataBanks_3_io_w_data_4),
    .io_w_data_5(dataBanks_3_io_w_data_5),
    .io_w_data_6(dataBanks_3_io_w_data_6),
    .io_w_data_7(dataBanks_3_io_w_data_7),
    .io_w_maskOH(dataBanks_3_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_4 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_4_clock),
    .reset(dataBanks_4_reset),
    .io_r_addr(dataBanks_4_io_r_addr),
    .io_r_data_0(dataBanks_4_io_r_data_0),
    .io_r_data_1(dataBanks_4_io_r_data_1),
    .io_r_data_2(dataBanks_4_io_r_data_2),
    .io_r_data_3(dataBanks_4_io_r_data_3),
    .io_r_data_4(dataBanks_4_io_r_data_4),
    .io_r_data_5(dataBanks_4_io_r_data_5),
    .io_r_data_6(dataBanks_4_io_r_data_6),
    .io_r_data_7(dataBanks_4_io_r_data_7),
    .io_w_en(dataBanks_4_io_w_en),
    .io_w_addr(dataBanks_4_io_w_addr),
    .io_w_data_0(dataBanks_4_io_w_data_0),
    .io_w_data_1(dataBanks_4_io_w_data_1),
    .io_w_data_2(dataBanks_4_io_w_data_2),
    .io_w_data_3(dataBanks_4_io_w_data_3),
    .io_w_data_4(dataBanks_4_io_w_data_4),
    .io_w_data_5(dataBanks_4_io_w_data_5),
    .io_w_data_6(dataBanks_4_io_w_data_6),
    .io_w_data_7(dataBanks_4_io_w_data_7),
    .io_w_maskOH(dataBanks_4_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_5 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_5_clock),
    .reset(dataBanks_5_reset),
    .io_r_addr(dataBanks_5_io_r_addr),
    .io_r_data_0(dataBanks_5_io_r_data_0),
    .io_r_data_1(dataBanks_5_io_r_data_1),
    .io_r_data_2(dataBanks_5_io_r_data_2),
    .io_r_data_3(dataBanks_5_io_r_data_3),
    .io_r_data_4(dataBanks_5_io_r_data_4),
    .io_r_data_5(dataBanks_5_io_r_data_5),
    .io_r_data_6(dataBanks_5_io_r_data_6),
    .io_r_data_7(dataBanks_5_io_r_data_7),
    .io_w_en(dataBanks_5_io_w_en),
    .io_w_addr(dataBanks_5_io_w_addr),
    .io_w_data_0(dataBanks_5_io_w_data_0),
    .io_w_data_1(dataBanks_5_io_w_data_1),
    .io_w_data_2(dataBanks_5_io_w_data_2),
    .io_w_data_3(dataBanks_5_io_w_data_3),
    .io_w_data_4(dataBanks_5_io_w_data_4),
    .io_w_data_5(dataBanks_5_io_w_data_5),
    .io_w_data_6(dataBanks_5_io_w_data_6),
    .io_w_data_7(dataBanks_5_io_w_data_7),
    .io_w_maskOH(dataBanks_5_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_6 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_6_clock),
    .reset(dataBanks_6_reset),
    .io_r_addr(dataBanks_6_io_r_addr),
    .io_r_data_0(dataBanks_6_io_r_data_0),
    .io_r_data_1(dataBanks_6_io_r_data_1),
    .io_r_data_2(dataBanks_6_io_r_data_2),
    .io_r_data_3(dataBanks_6_io_r_data_3),
    .io_r_data_4(dataBanks_6_io_r_data_4),
    .io_r_data_5(dataBanks_6_io_r_data_5),
    .io_r_data_6(dataBanks_6_io_r_data_6),
    .io_r_data_7(dataBanks_6_io_r_data_7),
    .io_w_en(dataBanks_6_io_w_en),
    .io_w_addr(dataBanks_6_io_w_addr),
    .io_w_data_0(dataBanks_6_io_w_data_0),
    .io_w_data_1(dataBanks_6_io_w_data_1),
    .io_w_data_2(dataBanks_6_io_w_data_2),
    .io_w_data_3(dataBanks_6_io_w_data_3),
    .io_w_data_4(dataBanks_6_io_w_data_4),
    .io_w_data_5(dataBanks_6_io_w_data_5),
    .io_w_data_6(dataBanks_6_io_w_data_6),
    .io_w_data_7(dataBanks_6_io_w_data_7),
    .io_w_maskOH(dataBanks_6_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_7 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_7_clock),
    .reset(dataBanks_7_reset),
    .io_r_addr(dataBanks_7_io_r_addr),
    .io_r_data_0(dataBanks_7_io_r_data_0),
    .io_r_data_1(dataBanks_7_io_r_data_1),
    .io_r_data_2(dataBanks_7_io_r_data_2),
    .io_r_data_3(dataBanks_7_io_r_data_3),
    .io_r_data_4(dataBanks_7_io_r_data_4),
    .io_r_data_5(dataBanks_7_io_r_data_5),
    .io_r_data_6(dataBanks_7_io_r_data_6),
    .io_r_data_7(dataBanks_7_io_r_data_7),
    .io_w_en(dataBanks_7_io_w_en),
    .io_w_addr(dataBanks_7_io_w_addr),
    .io_w_data_0(dataBanks_7_io_w_data_0),
    .io_w_data_1(dataBanks_7_io_w_data_1),
    .io_w_data_2(dataBanks_7_io_w_data_2),
    .io_w_data_3(dataBanks_7_io_w_data_3),
    .io_w_data_4(dataBanks_7_io_w_data_4),
    .io_w_data_5(dataBanks_7_io_w_data_5),
    .io_w_data_6(dataBanks_7_io_w_data_6),
    .io_w_data_7(dataBanks_7_io_w_data_7),
    .io_w_maskOH(dataBanks_7_io_w_maskOH)
  );
  assign io_read_req_ready = 1'h1; // @[DataBank.scala 46:23]
  assign io_read_resp_0_0 = ren ? dataBanks_0_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_1 = ren ? dataBanks_0_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_2 = ren ? dataBanks_0_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_3 = ren ? dataBanks_0_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_4 = ren ? dataBanks_0_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_5 = ren ? dataBanks_0_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_6 = ren ? dataBanks_0_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_7 = ren ? dataBanks_0_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_0 = ren ? dataBanks_1_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_1 = ren ? dataBanks_1_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_2 = ren ? dataBanks_1_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_3 = ren ? dataBanks_1_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_4 = ren ? dataBanks_1_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_5 = ren ? dataBanks_1_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_6 = ren ? dataBanks_1_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_7 = ren ? dataBanks_1_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_0 = ren ? dataBanks_2_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_1 = ren ? dataBanks_2_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_2 = ren ? dataBanks_2_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_3 = ren ? dataBanks_2_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_4 = ren ? dataBanks_2_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_5 = ren ? dataBanks_2_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_6 = ren ? dataBanks_2_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_7 = ren ? dataBanks_2_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_0 = ren ? dataBanks_3_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_1 = ren ? dataBanks_3_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_2 = ren ? dataBanks_3_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_3 = ren ? dataBanks_3_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_4 = ren ? dataBanks_3_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_5 = ren ? dataBanks_3_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_6 = ren ? dataBanks_3_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_7 = ren ? dataBanks_3_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_0 = ren ? dataBanks_4_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_1 = ren ? dataBanks_4_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_2 = ren ? dataBanks_4_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_3 = ren ? dataBanks_4_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_4 = ren ? dataBanks_4_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_5 = ren ? dataBanks_4_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_6 = ren ? dataBanks_4_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_7 = ren ? dataBanks_4_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_0 = ren ? dataBanks_5_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_1 = ren ? dataBanks_5_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_2 = ren ? dataBanks_5_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_3 = ren ? dataBanks_5_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_4 = ren ? dataBanks_5_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_5 = ren ? dataBanks_5_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_6 = ren ? dataBanks_5_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_7 = ren ? dataBanks_5_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_0 = ren ? dataBanks_6_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_1 = ren ? dataBanks_6_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_2 = ren ? dataBanks_6_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_3 = ren ? dataBanks_6_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_4 = ren ? dataBanks_6_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_5 = ren ? dataBanks_6_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_6 = ren ? dataBanks_6_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_7 = ren ? dataBanks_6_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_0 = ren ? dataBanks_7_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_1 = ren ? dataBanks_7_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_2 = ren ? dataBanks_7_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_3 = ren ? dataBanks_7_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_4 = ren ? dataBanks_7_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_5 = ren ? dataBanks_7_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_6 = ren ? dataBanks_7_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_7 = ren ? dataBanks_7_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_write_req_ready = 1'h1; // @[DataBank.scala 55:28]
  assign dataBanks_0_clock = clock;
  assign dataBanks_0_reset = reset;
  assign dataBanks_0_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_0_io_w_en = io_write_req_bits_way[0] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_0_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_0_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_1_clock = clock;
  assign dataBanks_1_reset = reset;
  assign dataBanks_1_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_1_io_w_en = io_write_req_bits_way[1] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_1_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_1_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_2_clock = clock;
  assign dataBanks_2_reset = reset;
  assign dataBanks_2_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_2_io_w_en = io_write_req_bits_way[2] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_2_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_2_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_3_clock = clock;
  assign dataBanks_3_reset = reset;
  assign dataBanks_3_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_3_io_w_en = io_write_req_bits_way[3] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_3_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_3_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_4_clock = clock;
  assign dataBanks_4_reset = reset;
  assign dataBanks_4_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_4_io_w_en = io_write_req_bits_way[4] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_4_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_4_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_5_clock = clock;
  assign dataBanks_5_reset = reset;
  assign dataBanks_5_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_5_io_w_en = io_write_req_bits_way[5] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_5_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_5_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_6_clock = clock;
  assign dataBanks_6_reset = reset;
  assign dataBanks_6_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_6_io_w_en = io_write_req_bits_way[6] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_6_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_6_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_7_clock = clock;
  assign dataBanks_7_reset = reset;
  assign dataBanks_7_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_7_io_w_en = io_write_req_bits_way[7] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_7_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_7_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
endmodule
module BankRAM_2P_64(
  input         clock,
  input         reset,
  input  [6:0]  io_r_addr,
  output [19:0] io_r_data,
  input         io_w_en,
  input  [6:0]  io_w_addr,
  input  [19:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] mem [0:127]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [6:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 20'h0;
  assign mem_MPORT_addr = 7'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 20'h0;
  assign mem_MPORT_1_addr = 7'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 20'h0;
  assign mem_MPORT_2_addr = 7'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 20'h0;
  assign mem_MPORT_3_addr = 7'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 20'h0;
  assign mem_MPORT_4_addr = 7'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 20'h0;
  assign mem_MPORT_5_addr = 7'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 20'h0;
  assign mem_MPORT_6_addr = 7'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 20'h0;
  assign mem_MPORT_7_addr = 7'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 20'h0;
  assign mem_MPORT_8_addr = 7'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 20'h0;
  assign mem_MPORT_9_addr = 7'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 20'h0;
  assign mem_MPORT_10_addr = 7'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 20'h0;
  assign mem_MPORT_11_addr = 7'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 20'h0;
  assign mem_MPORT_12_addr = 7'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 20'h0;
  assign mem_MPORT_13_addr = 7'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 20'h0;
  assign mem_MPORT_14_addr = 7'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 20'h0;
  assign mem_MPORT_15_addr = 7'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 20'h0;
  assign mem_MPORT_16_addr = 7'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 20'h0;
  assign mem_MPORT_17_addr = 7'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 20'h0;
  assign mem_MPORT_18_addr = 7'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 20'h0;
  assign mem_MPORT_19_addr = 7'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 20'h0;
  assign mem_MPORT_20_addr = 7'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 20'h0;
  assign mem_MPORT_21_addr = 7'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 20'h0;
  assign mem_MPORT_22_addr = 7'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 20'h0;
  assign mem_MPORT_23_addr = 7'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 20'h0;
  assign mem_MPORT_24_addr = 7'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 20'h0;
  assign mem_MPORT_25_addr = 7'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 20'h0;
  assign mem_MPORT_26_addr = 7'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 20'h0;
  assign mem_MPORT_27_addr = 7'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 20'h0;
  assign mem_MPORT_28_addr = 7'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 20'h0;
  assign mem_MPORT_29_addr = 7'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 20'h0;
  assign mem_MPORT_30_addr = 7'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 20'h0;
  assign mem_MPORT_31_addr = 7'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 20'h0;
  assign mem_MPORT_32_addr = 7'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 20'h0;
  assign mem_MPORT_33_addr = 7'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 20'h0;
  assign mem_MPORT_34_addr = 7'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 20'h0;
  assign mem_MPORT_35_addr = 7'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 20'h0;
  assign mem_MPORT_36_addr = 7'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 20'h0;
  assign mem_MPORT_37_addr = 7'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 20'h0;
  assign mem_MPORT_38_addr = 7'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 20'h0;
  assign mem_MPORT_39_addr = 7'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 20'h0;
  assign mem_MPORT_40_addr = 7'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 20'h0;
  assign mem_MPORT_41_addr = 7'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 20'h0;
  assign mem_MPORT_42_addr = 7'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 20'h0;
  assign mem_MPORT_43_addr = 7'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 20'h0;
  assign mem_MPORT_44_addr = 7'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 20'h0;
  assign mem_MPORT_45_addr = 7'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 20'h0;
  assign mem_MPORT_46_addr = 7'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 20'h0;
  assign mem_MPORT_47_addr = 7'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 20'h0;
  assign mem_MPORT_48_addr = 7'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 20'h0;
  assign mem_MPORT_49_addr = 7'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 20'h0;
  assign mem_MPORT_50_addr = 7'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 20'h0;
  assign mem_MPORT_51_addr = 7'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 20'h0;
  assign mem_MPORT_52_addr = 7'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 20'h0;
  assign mem_MPORT_53_addr = 7'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 20'h0;
  assign mem_MPORT_54_addr = 7'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 20'h0;
  assign mem_MPORT_55_addr = 7'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 20'h0;
  assign mem_MPORT_56_addr = 7'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 20'h0;
  assign mem_MPORT_57_addr = 7'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 20'h0;
  assign mem_MPORT_58_addr = 7'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 20'h0;
  assign mem_MPORT_59_addr = 7'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 20'h0;
  assign mem_MPORT_60_addr = 7'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 20'h0;
  assign mem_MPORT_61_addr = 7'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 20'h0;
  assign mem_MPORT_62_addr = 7'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 20'h0;
  assign mem_MPORT_63_addr = 7'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 20'h0;
  assign mem_MPORT_64_addr = 7'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 20'h0;
  assign mem_MPORT_65_addr = 7'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 20'h0;
  assign mem_MPORT_66_addr = 7'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 20'h0;
  assign mem_MPORT_67_addr = 7'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 20'h0;
  assign mem_MPORT_68_addr = 7'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 20'h0;
  assign mem_MPORT_69_addr = 7'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 20'h0;
  assign mem_MPORT_70_addr = 7'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 20'h0;
  assign mem_MPORT_71_addr = 7'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 20'h0;
  assign mem_MPORT_72_addr = 7'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 20'h0;
  assign mem_MPORT_73_addr = 7'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 20'h0;
  assign mem_MPORT_74_addr = 7'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 20'h0;
  assign mem_MPORT_75_addr = 7'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 20'h0;
  assign mem_MPORT_76_addr = 7'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 20'h0;
  assign mem_MPORT_77_addr = 7'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 20'h0;
  assign mem_MPORT_78_addr = 7'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 20'h0;
  assign mem_MPORT_79_addr = 7'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 20'h0;
  assign mem_MPORT_80_addr = 7'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 20'h0;
  assign mem_MPORT_81_addr = 7'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 20'h0;
  assign mem_MPORT_82_addr = 7'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 20'h0;
  assign mem_MPORT_83_addr = 7'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 20'h0;
  assign mem_MPORT_84_addr = 7'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 20'h0;
  assign mem_MPORT_85_addr = 7'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 20'h0;
  assign mem_MPORT_86_addr = 7'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 20'h0;
  assign mem_MPORT_87_addr = 7'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 20'h0;
  assign mem_MPORT_88_addr = 7'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 20'h0;
  assign mem_MPORT_89_addr = 7'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 20'h0;
  assign mem_MPORT_90_addr = 7'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 20'h0;
  assign mem_MPORT_91_addr = 7'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 20'h0;
  assign mem_MPORT_92_addr = 7'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 20'h0;
  assign mem_MPORT_93_addr = 7'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 20'h0;
  assign mem_MPORT_94_addr = 7'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 20'h0;
  assign mem_MPORT_95_addr = 7'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 20'h0;
  assign mem_MPORT_96_addr = 7'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 20'h0;
  assign mem_MPORT_97_addr = 7'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 20'h0;
  assign mem_MPORT_98_addr = 7'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 20'h0;
  assign mem_MPORT_99_addr = 7'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 20'h0;
  assign mem_MPORT_100_addr = 7'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 20'h0;
  assign mem_MPORT_101_addr = 7'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 20'h0;
  assign mem_MPORT_102_addr = 7'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 20'h0;
  assign mem_MPORT_103_addr = 7'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 20'h0;
  assign mem_MPORT_104_addr = 7'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 20'h0;
  assign mem_MPORT_105_addr = 7'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 20'h0;
  assign mem_MPORT_106_addr = 7'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 20'h0;
  assign mem_MPORT_107_addr = 7'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 20'h0;
  assign mem_MPORT_108_addr = 7'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 20'h0;
  assign mem_MPORT_109_addr = 7'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 20'h0;
  assign mem_MPORT_110_addr = 7'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 20'h0;
  assign mem_MPORT_111_addr = 7'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 20'h0;
  assign mem_MPORT_112_addr = 7'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 20'h0;
  assign mem_MPORT_113_addr = 7'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 20'h0;
  assign mem_MPORT_114_addr = 7'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 20'h0;
  assign mem_MPORT_115_addr = 7'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 20'h0;
  assign mem_MPORT_116_addr = 7'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 20'h0;
  assign mem_MPORT_117_addr = 7'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 20'h0;
  assign mem_MPORT_118_addr = 7'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 20'h0;
  assign mem_MPORT_119_addr = 7'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 20'h0;
  assign mem_MPORT_120_addr = 7'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 20'h0;
  assign mem_MPORT_121_addr = 7'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 20'h0;
  assign mem_MPORT_122_addr = 7'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 20'h0;
  assign mem_MPORT_123_addr = 7'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 20'h0;
  assign mem_MPORT_124_addr = 7'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 20'h0;
  assign mem_MPORT_125_addr = 7'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 20'h0;
  assign mem_MPORT_126_addr = 7'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 20'h0;
  assign mem_MPORT_127_addr = 7'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = io_w_data;
  assign mem_MPORT_128_addr = io_w_addr;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_8(
  input         clock,
  input         reset,
  input  [6:0]  io_r_addr,
  output [19:0] io_r_data_0,
  output [19:0] io_r_data_1,
  output [19:0] io_r_data_2,
  output [19:0] io_r_data_3,
  output [19:0] io_r_data_4,
  output [19:0] io_r_data_5,
  output [19:0] io_r_data_6,
  output [19:0] io_r_data_7,
  input         io_w_en,
  input  [6:0]  io_w_addr,
  input  [19:0] io_w_data_0,
  input  [19:0] io_w_data_1,
  input  [19:0] io_w_data_2,
  input  [19:0] io_w_data_3,
  input  [19:0] io_w_data_4,
  input  [19:0] io_w_data_5,
  input  [19:0] io_w_data_6,
  input  [19:0] io_w_data_7,
  input  [7:0]  io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_clock; // @[SRAM_1.scala 201:38]
  wire  brams_4_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_4_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_4_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_clock; // @[SRAM_1.scala 201:38]
  wire  brams_5_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_5_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_5_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_clock; // @[SRAM_1.scala 201:38]
  wire  brams_6_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_6_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_6_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_clock; // @[SRAM_1.scala 201:38]
  wire  brams_7_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_7_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_7_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P_64 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P_64 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P_64 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P_64 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  BankRAM_2P_64 brams_4 ( // @[SRAM_1.scala 201:38]
    .clock(brams_4_clock),
    .reset(brams_4_reset),
    .io_r_addr(brams_4_io_r_addr),
    .io_r_data(brams_4_io_r_data),
    .io_w_en(brams_4_io_w_en),
    .io_w_addr(brams_4_io_w_addr),
    .io_w_data(brams_4_io_w_data)
  );
  BankRAM_2P_64 brams_5 ( // @[SRAM_1.scala 201:38]
    .clock(brams_5_clock),
    .reset(brams_5_reset),
    .io_r_addr(brams_5_io_r_addr),
    .io_r_data(brams_5_io_r_data),
    .io_w_en(brams_5_io_w_en),
    .io_w_addr(brams_5_io_w_addr),
    .io_w_data(brams_5_io_w_data)
  );
  BankRAM_2P_64 brams_6 ( // @[SRAM_1.scala 201:38]
    .clock(brams_6_clock),
    .reset(brams_6_reset),
    .io_r_addr(brams_6_io_r_addr),
    .io_r_data(brams_6_io_r_data),
    .io_w_en(brams_6_io_w_en),
    .io_w_addr(brams_6_io_w_addr),
    .io_w_data(brams_6_io_w_data)
  );
  BankRAM_2P_64 brams_7 ( // @[SRAM_1.scala 201:38]
    .clock(brams_7_clock),
    .reset(brams_7_reset),
    .io_r_addr(brams_7_io_r_addr),
    .io_r_data(brams_7_io_r_data),
    .io_w_en(brams_7_io_w_en),
    .io_w_addr(brams_7_io_w_addr),
    .io_w_data(brams_7_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_4 = brams_4_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_5 = brams_5_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_6 = brams_6_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_7 = brams_7_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
  assign brams_4_clock = clock;
  assign brams_4_reset = reset;
  assign brams_4_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_4_io_w_en = io_w_en & io_w_maskOH[4]; // @[SRAM_1.scala 208:37]
  assign brams_4_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_4_io_w_data = io_w_data_4; // @[SRAM_1.scala 210:28]
  assign brams_5_clock = clock;
  assign brams_5_reset = reset;
  assign brams_5_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_5_io_w_en = io_w_en & io_w_maskOH[5]; // @[SRAM_1.scala 208:37]
  assign brams_5_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_5_io_w_data = io_w_data_5; // @[SRAM_1.scala 210:28]
  assign brams_6_clock = clock;
  assign brams_6_reset = reset;
  assign brams_6_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_6_io_w_en = io_w_en & io_w_maskOH[6]; // @[SRAM_1.scala 208:37]
  assign brams_6_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_6_io_w_data = io_w_data_6; // @[SRAM_1.scala 210:28]
  assign brams_7_clock = clock;
  assign brams_7_reset = reset;
  assign brams_7_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_7_io_w_en = io_w_en & io_w_maskOH[7]; // @[SRAM_1.scala 208:37]
  assign brams_7_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_7_io_w_data = io_w_data_7; // @[SRAM_1.scala 210:28]
endmodule
module BankRAM_2P_72(
  input        clock,
  input        reset,
  input  [6:0] io_r_addr,
  output [1:0] io_r_data,
  input        io_w_en,
  input  [6:0] io_w_addr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] mem [0:127]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [6:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 2'h0;
  assign mem_MPORT_addr = 7'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 2'h0;
  assign mem_MPORT_1_addr = 7'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 2'h0;
  assign mem_MPORT_2_addr = 7'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 2'h0;
  assign mem_MPORT_3_addr = 7'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 2'h0;
  assign mem_MPORT_4_addr = 7'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 2'h0;
  assign mem_MPORT_5_addr = 7'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 2'h0;
  assign mem_MPORT_6_addr = 7'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 2'h0;
  assign mem_MPORT_7_addr = 7'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 2'h0;
  assign mem_MPORT_8_addr = 7'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 2'h0;
  assign mem_MPORT_9_addr = 7'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 2'h0;
  assign mem_MPORT_10_addr = 7'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 2'h0;
  assign mem_MPORT_11_addr = 7'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 2'h0;
  assign mem_MPORT_12_addr = 7'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 2'h0;
  assign mem_MPORT_13_addr = 7'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 2'h0;
  assign mem_MPORT_14_addr = 7'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 2'h0;
  assign mem_MPORT_15_addr = 7'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 2'h0;
  assign mem_MPORT_16_addr = 7'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 2'h0;
  assign mem_MPORT_17_addr = 7'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 2'h0;
  assign mem_MPORT_18_addr = 7'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 2'h0;
  assign mem_MPORT_19_addr = 7'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 2'h0;
  assign mem_MPORT_20_addr = 7'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 2'h0;
  assign mem_MPORT_21_addr = 7'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 2'h0;
  assign mem_MPORT_22_addr = 7'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 2'h0;
  assign mem_MPORT_23_addr = 7'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 2'h0;
  assign mem_MPORT_24_addr = 7'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 2'h0;
  assign mem_MPORT_25_addr = 7'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 2'h0;
  assign mem_MPORT_26_addr = 7'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 2'h0;
  assign mem_MPORT_27_addr = 7'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 2'h0;
  assign mem_MPORT_28_addr = 7'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 2'h0;
  assign mem_MPORT_29_addr = 7'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 2'h0;
  assign mem_MPORT_30_addr = 7'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 2'h0;
  assign mem_MPORT_31_addr = 7'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 2'h0;
  assign mem_MPORT_32_addr = 7'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 2'h0;
  assign mem_MPORT_33_addr = 7'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 2'h0;
  assign mem_MPORT_34_addr = 7'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 2'h0;
  assign mem_MPORT_35_addr = 7'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 2'h0;
  assign mem_MPORT_36_addr = 7'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 2'h0;
  assign mem_MPORT_37_addr = 7'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 2'h0;
  assign mem_MPORT_38_addr = 7'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 2'h0;
  assign mem_MPORT_39_addr = 7'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 2'h0;
  assign mem_MPORT_40_addr = 7'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 2'h0;
  assign mem_MPORT_41_addr = 7'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 2'h0;
  assign mem_MPORT_42_addr = 7'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 2'h0;
  assign mem_MPORT_43_addr = 7'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 2'h0;
  assign mem_MPORT_44_addr = 7'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 2'h0;
  assign mem_MPORT_45_addr = 7'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 2'h0;
  assign mem_MPORT_46_addr = 7'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 2'h0;
  assign mem_MPORT_47_addr = 7'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 2'h0;
  assign mem_MPORT_48_addr = 7'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 2'h0;
  assign mem_MPORT_49_addr = 7'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 2'h0;
  assign mem_MPORT_50_addr = 7'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 2'h0;
  assign mem_MPORT_51_addr = 7'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 2'h0;
  assign mem_MPORT_52_addr = 7'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 2'h0;
  assign mem_MPORT_53_addr = 7'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 2'h0;
  assign mem_MPORT_54_addr = 7'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 2'h0;
  assign mem_MPORT_55_addr = 7'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 2'h0;
  assign mem_MPORT_56_addr = 7'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 2'h0;
  assign mem_MPORT_57_addr = 7'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 2'h0;
  assign mem_MPORT_58_addr = 7'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 2'h0;
  assign mem_MPORT_59_addr = 7'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 2'h0;
  assign mem_MPORT_60_addr = 7'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 2'h0;
  assign mem_MPORT_61_addr = 7'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 2'h0;
  assign mem_MPORT_62_addr = 7'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 2'h0;
  assign mem_MPORT_63_addr = 7'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 2'h0;
  assign mem_MPORT_64_addr = 7'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 2'h0;
  assign mem_MPORT_65_addr = 7'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 2'h0;
  assign mem_MPORT_66_addr = 7'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 2'h0;
  assign mem_MPORT_67_addr = 7'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 2'h0;
  assign mem_MPORT_68_addr = 7'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 2'h0;
  assign mem_MPORT_69_addr = 7'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 2'h0;
  assign mem_MPORT_70_addr = 7'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 2'h0;
  assign mem_MPORT_71_addr = 7'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 2'h0;
  assign mem_MPORT_72_addr = 7'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 2'h0;
  assign mem_MPORT_73_addr = 7'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 2'h0;
  assign mem_MPORT_74_addr = 7'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 2'h0;
  assign mem_MPORT_75_addr = 7'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 2'h0;
  assign mem_MPORT_76_addr = 7'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 2'h0;
  assign mem_MPORT_77_addr = 7'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 2'h0;
  assign mem_MPORT_78_addr = 7'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 2'h0;
  assign mem_MPORT_79_addr = 7'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 2'h0;
  assign mem_MPORT_80_addr = 7'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 2'h0;
  assign mem_MPORT_81_addr = 7'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 2'h0;
  assign mem_MPORT_82_addr = 7'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 2'h0;
  assign mem_MPORT_83_addr = 7'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 2'h0;
  assign mem_MPORT_84_addr = 7'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 2'h0;
  assign mem_MPORT_85_addr = 7'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 2'h0;
  assign mem_MPORT_86_addr = 7'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 2'h0;
  assign mem_MPORT_87_addr = 7'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 2'h0;
  assign mem_MPORT_88_addr = 7'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 2'h0;
  assign mem_MPORT_89_addr = 7'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 2'h0;
  assign mem_MPORT_90_addr = 7'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 2'h0;
  assign mem_MPORT_91_addr = 7'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 2'h0;
  assign mem_MPORT_92_addr = 7'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 2'h0;
  assign mem_MPORT_93_addr = 7'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 2'h0;
  assign mem_MPORT_94_addr = 7'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 2'h0;
  assign mem_MPORT_95_addr = 7'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 2'h0;
  assign mem_MPORT_96_addr = 7'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 2'h0;
  assign mem_MPORT_97_addr = 7'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 2'h0;
  assign mem_MPORT_98_addr = 7'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 2'h0;
  assign mem_MPORT_99_addr = 7'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 2'h0;
  assign mem_MPORT_100_addr = 7'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 2'h0;
  assign mem_MPORT_101_addr = 7'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 2'h0;
  assign mem_MPORT_102_addr = 7'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 2'h0;
  assign mem_MPORT_103_addr = 7'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 2'h0;
  assign mem_MPORT_104_addr = 7'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 2'h0;
  assign mem_MPORT_105_addr = 7'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 2'h0;
  assign mem_MPORT_106_addr = 7'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 2'h0;
  assign mem_MPORT_107_addr = 7'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 2'h0;
  assign mem_MPORT_108_addr = 7'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 2'h0;
  assign mem_MPORT_109_addr = 7'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 2'h0;
  assign mem_MPORT_110_addr = 7'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 2'h0;
  assign mem_MPORT_111_addr = 7'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 2'h0;
  assign mem_MPORT_112_addr = 7'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 2'h0;
  assign mem_MPORT_113_addr = 7'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 2'h0;
  assign mem_MPORT_114_addr = 7'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 2'h0;
  assign mem_MPORT_115_addr = 7'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 2'h0;
  assign mem_MPORT_116_addr = 7'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 2'h0;
  assign mem_MPORT_117_addr = 7'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 2'h0;
  assign mem_MPORT_118_addr = 7'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 2'h0;
  assign mem_MPORT_119_addr = 7'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 2'h0;
  assign mem_MPORT_120_addr = 7'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 2'h0;
  assign mem_MPORT_121_addr = 7'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 2'h0;
  assign mem_MPORT_122_addr = 7'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 2'h0;
  assign mem_MPORT_123_addr = 7'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 2'h0;
  assign mem_MPORT_124_addr = 7'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 2'h0;
  assign mem_MPORT_125_addr = 7'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 2'h0;
  assign mem_MPORT_126_addr = 7'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 2'h0;
  assign mem_MPORT_127_addr = 7'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 2'h1;
  assign mem_MPORT_128_addr = io_w_addr;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? 2'h1 : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_9(
  input        clock,
  input        reset,
  input  [6:0] io_r_addr,
  output [1:0] io_r_data_0,
  output [1:0] io_r_data_1,
  output [1:0] io_r_data_2,
  output [1:0] io_r_data_3,
  output [1:0] io_r_data_4,
  output [1:0] io_r_data_5,
  output [1:0] io_r_data_6,
  output [1:0] io_r_data_7,
  input        io_w_en,
  input  [6:0] io_w_addr,
  input  [7:0] io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_4_clock; // @[SRAM_1.scala 201:38]
  wire  brams_4_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_4_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_5_clock; // @[SRAM_1.scala 201:38]
  wire  brams_5_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_5_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_6_clock; // @[SRAM_1.scala 201:38]
  wire  brams_6_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_6_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_7_clock; // @[SRAM_1.scala 201:38]
  wire  brams_7_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_7_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_w_addr; // @[SRAM_1.scala 201:38]
  BankRAM_2P_72 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr)
  );
  BankRAM_2P_72 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr)
  );
  BankRAM_2P_72 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr)
  );
  BankRAM_2P_72 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr)
  );
  BankRAM_2P_72 brams_4 ( // @[SRAM_1.scala 201:38]
    .clock(brams_4_clock),
    .reset(brams_4_reset),
    .io_r_addr(brams_4_io_r_addr),
    .io_r_data(brams_4_io_r_data),
    .io_w_en(brams_4_io_w_en),
    .io_w_addr(brams_4_io_w_addr)
  );
  BankRAM_2P_72 brams_5 ( // @[SRAM_1.scala 201:38]
    .clock(brams_5_clock),
    .reset(brams_5_reset),
    .io_r_addr(brams_5_io_r_addr),
    .io_r_data(brams_5_io_r_data),
    .io_w_en(brams_5_io_w_en),
    .io_w_addr(brams_5_io_w_addr)
  );
  BankRAM_2P_72 brams_6 ( // @[SRAM_1.scala 201:38]
    .clock(brams_6_clock),
    .reset(brams_6_reset),
    .io_r_addr(brams_6_io_r_addr),
    .io_r_data(brams_6_io_r_data),
    .io_w_en(brams_6_io_w_en),
    .io_w_addr(brams_6_io_w_addr)
  );
  BankRAM_2P_72 brams_7 ( // @[SRAM_1.scala 201:38]
    .clock(brams_7_clock),
    .reset(brams_7_reset),
    .io_r_addr(brams_7_io_r_addr),
    .io_r_data(brams_7_io_r_data),
    .io_w_en(brams_7_io_w_en),
    .io_w_addr(brams_7_io_w_addr)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_4 = brams_4_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_5 = brams_5_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_6 = brams_6_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_7 = brams_7_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_4_clock = clock;
  assign brams_4_reset = reset;
  assign brams_4_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_4_io_w_en = io_w_en & io_w_maskOH[4]; // @[SRAM_1.scala 208:37]
  assign brams_4_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_5_clock = clock;
  assign brams_5_reset = reset;
  assign brams_5_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_5_io_w_en = io_w_en & io_w_maskOH[5]; // @[SRAM_1.scala 208:37]
  assign brams_5_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_6_clock = clock;
  assign brams_6_reset = reset;
  assign brams_6_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_6_io_w_en = io_w_en & io_w_maskOH[6]; // @[SRAM_1.scala 208:37]
  assign brams_6_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_7_clock = clock;
  assign brams_7_reset = reset;
  assign brams_7_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_7_io_w_en = io_w_en & io_w_maskOH[7]; // @[SRAM_1.scala 208:37]
  assign brams_7_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  reg  state_8; // @[PRNG.scala 55:49]
  reg  state_9; // @[PRNG.scala 55:49]
  reg  state_10; // @[PRNG.scala 55:49]
  reg  state_11; // @[PRNG.scala 55:49]
  reg  state_12; // @[PRNG.scala 55:49]
  reg  state_13; // @[PRNG.scala 55:49]
  reg  state_14; // @[PRNG.scala 55:49]
  reg  state_15; // @[PRNG.scala 55:49]
  wire  _T_2 = state_15 ^ state_13 ^ state_12 ^ state_10; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  assign io_out_8 = state_8; // @[PRNG.scala 78:10]
  assign io_out_9 = state_9; // @[PRNG.scala 78:10]
  assign io_out_10 = state_10; // @[PRNG.scala 78:10]
  assign io_out_11 = state_11; // @[PRNG.scala 78:10]
  assign io_out_12 = state_12; // @[PRNG.scala 78:10]
  assign io_out_13 = state_13; // @[PRNG.scala 78:10]
  assign io_out_14 = state_14; // @[PRNG.scala 78:10]
  assign io_out_15 = state_15; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T_2; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_4 <= state_3;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_5 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_5 <= state_4;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_6 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_6 <= state_5;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_7 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_7 <= state_6;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_8 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_8 <= state_7;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_9 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_9 <= state_8;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_10 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_10 <= state_9;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_11 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_11 <= state_10;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_12 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_12 <= state_11;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_13 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_13 <= state_12;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_14 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_14 <= state_13;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_15 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_15 <= state_14;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCacheDirectory(
  input         clock,
  input         reset,
  output        io_read_req_ready,
  input         io_read_req_valid,
  input  [31:0] io_read_req_bits_addr,
  output        io_read_resp_bits_hit,
  output [7:0]  io_read_resp_bits_chosenWay,
  output        io_write_req_ready,
  input         io_write_req_valid,
  input  [31:0] io_write_req_bits_addr,
  input  [7:0]  io_write_req_bits_way
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  tagArray_clock; // @[SRAM_1.scala 255:31]
  wire  tagArray_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] tagArray_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  tagArray_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] tagArray_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] tagArray_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  metaArray_clock; // @[SRAM_1.scala 255:31]
  wire  metaArray_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] metaArray_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  metaArray_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] metaArray_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [7:0] metaArray_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  replaceWay_lfsr_prng_clock; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_reset; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_15; // @[PRNG.scala 91:22]
  wire [6:0] rSet = io_read_req_bits_addr[11:5]; // @[Parameters.scala 50:11]
  wire [19:0] rTag = io_read_req_bits_addr[31:12]; // @[Parameters.scala 46:11]
  wire  ren = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  wire [6:0] wSet = io_write_req_bits_addr[11:5]; // @[Parameters.scala 50:11]
  wire [19:0] wTag = io_write_req_bits_addr[31:12]; // @[Parameters.scala 46:11]
  wire  wen = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _T_8 = io_write_req_bits_way[0] + io_write_req_bits_way[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_10 = io_write_req_bits_way[2] + io_write_req_bits_way[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_12 = _T_8 + _T_10; // @[Bitwise.scala 51:90]
  wire [1:0] _T_14 = io_write_req_bits_way[4] + io_write_req_bits_way[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_16 = io_write_req_bits_way[6] + io_write_req_bits_way[7]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_18 = _T_14 + _T_16; // @[Bitwise.scala 51:90]
  wire [3:0] _T_20 = _T_12 + _T_18; // @[Bitwise.scala 51:90]
  wire  _T_46 = ~reset; // @[Directory.scala 69:11]
  wire [19:0] rdata__0 = ren ? tagArray_io_r_data_0 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__1 = ren ? tagArray_io_r_data_1 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__2 = ren ? tagArray_io_r_data_2 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__3 = ren ? tagArray_io_r_data_3 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__4 = ren ? tagArray_io_r_data_4 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__5 = ren ? tagArray_io_r_data_5 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__6 = ren ? tagArray_io_r_data_6 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__7 = ren ? tagArray_io_r_data_7 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_0 = ren ? metaArray_io_r_data_0 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_1 = ren ? metaArray_io_r_data_1 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_2 = ren ? metaArray_io_r_data_2 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_3 = ren ? metaArray_io_r_data_3 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_4 = ren ? metaArray_io_r_data_4 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_5 = ren ? metaArray_io_r_data_5 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_6 = ren ? metaArray_io_r_data_6 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_7 = ren ? metaArray_io_r_data_7 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [15:0] _T_48 = {rdata_1_7,rdata_1_6,rdata_1_5,rdata_1_4,rdata_1_3,rdata_1_2,rdata_1_1,rdata_1_0}; // @[Directory.scala 82:52]
  wire  metaRdVec_0_valid = _T_48[0]; // @[Directory.scala 82:52]
  wire  metaRdVec_1_valid = _T_48[2]; // @[Directory.scala 82:52]
  wire  metaRdVec_2_valid = _T_48[4]; // @[Directory.scala 82:52]
  wire  metaRdVec_3_valid = _T_48[6]; // @[Directory.scala 82:52]
  wire  metaRdVec_4_valid = _T_48[8]; // @[Directory.scala 82:52]
  wire  metaRdVec_5_valid = _T_48[10]; // @[Directory.scala 82:52]
  wire  metaRdVec_6_valid = _T_48[12]; // @[Directory.scala 82:52]
  wire  metaRdVec_7_valid = _T_48[14]; // @[Directory.scala 82:52]
  wire  tagMatchVec_0 = rdata__0 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_1 = rdata__1 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_2 = rdata__2 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_3 = rdata__3 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_4 = rdata__4 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_5 = rdata__5 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_6 = rdata__6 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_7 = rdata__7 == rTag; // @[Directory.scala 85:46]
  wire  _matchWayOH_T = tagMatchVec_0 & metaRdVec_0_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_1 = tagMatchVec_1 & metaRdVec_1_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_2 = tagMatchVec_2 & metaRdVec_2_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_3 = tagMatchVec_3 & metaRdVec_3_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_4 = tagMatchVec_4 & metaRdVec_4_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_5 = tagMatchVec_5 & metaRdVec_5_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_6 = tagMatchVec_6 & metaRdVec_6_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_7 = tagMatchVec_7 & metaRdVec_7_valid; // @[Directory.scala 88:80]
  wire [7:0] matchWayOH = {_matchWayOH_T_7,_matchWayOH_T_6,_matchWayOH_T_5,_matchWayOH_T_4,_matchWayOH_T_3,
    _matchWayOH_T_2,_matchWayOH_T_1,_matchWayOH_T}; // @[Cat.scala 33:92]
  wire  invalidWayVec_0 = ~metaRdVec_0_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_1 = ~metaRdVec_1_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_2 = ~metaRdVec_2_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_3 = ~metaRdVec_3_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_4 = ~metaRdVec_4_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_5 = ~metaRdVec_5_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_6 = ~metaRdVec_6_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_7 = ~metaRdVec_7_valid; // @[Directory.scala 89:53]
  wire [7:0] _invalidWayOH_T_16 = invalidWayVec_6 ? 8'h40 : 8'h80; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_17 = invalidWayVec_5 ? 8'h20 : _invalidWayOH_T_16; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_18 = invalidWayVec_4 ? 8'h10 : _invalidWayOH_T_17; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_19 = invalidWayVec_3 ? 8'h8 : _invalidWayOH_T_18; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_20 = invalidWayVec_2 ? 8'h4 : _invalidWayOH_T_19; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_21 = invalidWayVec_1 ? 8'h2 : _invalidWayOH_T_20; // @[Mux.scala 47:70]
  wire [7:0] invalidWayOH = invalidWayVec_0 ? 8'h1 : _invalidWayOH_T_21; // @[Mux.scala 47:70]
  wire [7:0] _hasInvalidWay_T = {invalidWayVec_0,invalidWayVec_1,invalidWayVec_2,invalidWayVec_3,invalidWayVec_4,
    invalidWayVec_5,invalidWayVec_6,invalidWayVec_7}; // @[Cat.scala 33:92]
  wire  hasInvalidWay = |_hasInvalidWay_T; // @[Directory.scala 91:44]
  wire [7:0] replaceWay_lfsr_lo = {replaceWay_lfsr_prng_io_out_7,replaceWay_lfsr_prng_io_out_6,
    replaceWay_lfsr_prng_io_out_5,replaceWay_lfsr_prng_io_out_4,replaceWay_lfsr_prng_io_out_3,
    replaceWay_lfsr_prng_io_out_2,replaceWay_lfsr_prng_io_out_1,replaceWay_lfsr_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [15:0] replaceWay_lfsr = {replaceWay_lfsr_prng_io_out_15,replaceWay_lfsr_prng_io_out_14,
    replaceWay_lfsr_prng_io_out_13,replaceWay_lfsr_prng_io_out_12,replaceWay_lfsr_prng_io_out_11,
    replaceWay_lfsr_prng_io_out_10,replaceWay_lfsr_prng_io_out_9,replaceWay_lfsr_prng_io_out_8,replaceWay_lfsr_lo}; // @[PRNG.scala 95:17]
  wire [2:0] replaceWay_outputWay_shiftAmount = replaceWay_lfsr[2:0]; // @[DCache.scala 61:39]
  wire [7:0] replaceWay = 8'h1 << replaceWay_outputWay_shiftAmount; // @[OneHot.scala 64:12]
  wire  _replaceWayReg_T = ~io_read_req_valid; // @[Directory.scala 93:65]
  reg [7:0] replaceWayReg; // @[Reg.scala 19:16]
  wire  isHit = |matchWayOH; // @[Directory.scala 95:41]
  wire [7:0] _choseWayOH_T = hasInvalidWay ? invalidWayOH : replaceWayReg; // @[Directory.scala 96:51]
  wire [7:0] choseWayOH = isHit ? matchWayOH : _choseWayOH_T; // @[Directory.scala 96:28]
  wire [1:0] _T_73 = choseWayOH[0] + choseWayOH[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_75 = choseWayOH[2] + choseWayOH[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_77 = _T_73 + _T_75; // @[Bitwise.scala 51:90]
  wire [1:0] _T_79 = choseWayOH[4] + choseWayOH[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_81 = choseWayOH[6] + choseWayOH[7]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_83 = _T_79 + _T_81; // @[Bitwise.scala 51:90]
  wire [3:0] _T_85 = _T_77 + _T_83; // @[Bitwise.scala 51:90]
  SRAMArray_2P_8 tagArray ( // @[SRAM_1.scala 255:31]
    .clock(tagArray_clock),
    .reset(tagArray_reset),
    .io_r_addr(tagArray_io_r_addr),
    .io_r_data_0(tagArray_io_r_data_0),
    .io_r_data_1(tagArray_io_r_data_1),
    .io_r_data_2(tagArray_io_r_data_2),
    .io_r_data_3(tagArray_io_r_data_3),
    .io_r_data_4(tagArray_io_r_data_4),
    .io_r_data_5(tagArray_io_r_data_5),
    .io_r_data_6(tagArray_io_r_data_6),
    .io_r_data_7(tagArray_io_r_data_7),
    .io_w_en(tagArray_io_w_en),
    .io_w_addr(tagArray_io_w_addr),
    .io_w_data_0(tagArray_io_w_data_0),
    .io_w_data_1(tagArray_io_w_data_1),
    .io_w_data_2(tagArray_io_w_data_2),
    .io_w_data_3(tagArray_io_w_data_3),
    .io_w_data_4(tagArray_io_w_data_4),
    .io_w_data_5(tagArray_io_w_data_5),
    .io_w_data_6(tagArray_io_w_data_6),
    .io_w_data_7(tagArray_io_w_data_7),
    .io_w_maskOH(tagArray_io_w_maskOH)
  );
  SRAMArray_2P_9 metaArray ( // @[SRAM_1.scala 255:31]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_addr(metaArray_io_r_addr),
    .io_r_data_0(metaArray_io_r_data_0),
    .io_r_data_1(metaArray_io_r_data_1),
    .io_r_data_2(metaArray_io_r_data_2),
    .io_r_data_3(metaArray_io_r_data_3),
    .io_r_data_4(metaArray_io_r_data_4),
    .io_r_data_5(metaArray_io_r_data_5),
    .io_r_data_6(metaArray_io_r_data_6),
    .io_r_data_7(metaArray_io_r_data_7),
    .io_w_en(metaArray_io_w_en),
    .io_w_addr(metaArray_io_w_addr),
    .io_w_maskOH(metaArray_io_w_maskOH)
  );
  MaxPeriodFibonacciLFSR replaceWay_lfsr_prng ( // @[PRNG.scala 91:22]
    .clock(replaceWay_lfsr_prng_clock),
    .reset(replaceWay_lfsr_prng_reset),
    .io_out_0(replaceWay_lfsr_prng_io_out_0),
    .io_out_1(replaceWay_lfsr_prng_io_out_1),
    .io_out_2(replaceWay_lfsr_prng_io_out_2),
    .io_out_3(replaceWay_lfsr_prng_io_out_3),
    .io_out_4(replaceWay_lfsr_prng_io_out_4),
    .io_out_5(replaceWay_lfsr_prng_io_out_5),
    .io_out_6(replaceWay_lfsr_prng_io_out_6),
    .io_out_7(replaceWay_lfsr_prng_io_out_7),
    .io_out_8(replaceWay_lfsr_prng_io_out_8),
    .io_out_9(replaceWay_lfsr_prng_io_out_9),
    .io_out_10(replaceWay_lfsr_prng_io_out_10),
    .io_out_11(replaceWay_lfsr_prng_io_out_11),
    .io_out_12(replaceWay_lfsr_prng_io_out_12),
    .io_out_13(replaceWay_lfsr_prng_io_out_13),
    .io_out_14(replaceWay_lfsr_prng_io_out_14),
    .io_out_15(replaceWay_lfsr_prng_io_out_15)
  );
  assign io_read_req_ready = 1'h1; // @[Directory.scala 75:29]
  assign io_read_resp_bits_hit = |matchWayOH; // @[Directory.scala 95:41]
  assign io_read_resp_bits_chosenWay = isHit ? matchWayOH : _choseWayOH_T; // @[Directory.scala 96:28]
  assign io_write_req_ready = 1'h1; // @[Directory.scala 76:29]
  assign tagArray_clock = clock;
  assign tagArray_reset = reset;
  assign tagArray_io_r_addr = rSet; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign tagArray_io_w_en = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  assign tagArray_io_w_addr = wSet; // @[Directory.scala 112:15 SRAM_1.scala 237:19]
  assign tagArray_io_w_data_0 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_1 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_2 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_3 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_4 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_5 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_6 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_7 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_maskOH = io_write_req_bits_way; // @[Directory.scala 112:15 SRAM_1.scala 239:21]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r_addr = rSet; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign metaArray_io_w_en = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  assign metaArray_io_w_addr = wSet; // @[Directory.scala 112:15 SRAM_1.scala 237:19]
  assign metaArray_io_w_maskOH = io_write_req_bits_way; // @[Directory.scala 112:15 SRAM_1.scala 239:21]
  assign replaceWay_lfsr_prng_clock = clock;
  assign replaceWay_lfsr_prng_reset = reset;
  always @(posedge clock) begin
    if (_replaceWayReg_T) begin // @[Reg.scala 20:18]
      replaceWayReg <= replaceWay; // @[Reg.scala 20:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_20 < 4'h2)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Error directory write way has multiple valid bit! ==>%d\n    at Directory.scala:69 assert(PopCount(wWay) < 2.U, cf\"Error directory write way has multiple valid bit! ==>${PopCount(wWay)}\")\n"
            ,_T_20); // @[Directory.scala 69:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_20 < 4'h2) & ~reset) begin
          $fatal; // @[Directory.scala 69:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_46 & ~(_T_85 == 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Error chosenWay has multiple valid bit!\n    at Directory.scala:101 assert(PopCount(choseWayOH) === 1.U, \"Error chosenWay has multiple valid bit!\")\n"
            ); // @[Directory.scala 101:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_85 == 4'h1) & _T_46) begin
          $fatal; // @[Directory.scala 101:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wen & _T_46 & ~(_T_20 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: write error, tring to write multiple ways\n    at SRAM_1.scala:235 assert(PopCount(mask) <= 1.U, \"write error, tring to write multiple ways\")\n"
            ); // @[SRAM_1.scala 235:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_20 <= 4'h1) & (wen & _T_46)) begin
          $fatal; // @[SRAM_1.scala 235:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wen & _T_46 & ~(_T_20 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: write error, tring to write multiple ways\n    at SRAM_1.scala:235 assert(PopCount(mask) <= 1.U, \"write error, tring to write multiple ways\")\n"
            ); // @[SRAM_1.scala 235:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_20 <= 4'h1) & (wen & _T_46)) begin
          $fatal; // @[SRAM_1.scala 235:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  replaceWayReg = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RefillPipe(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [31:0]  io_req_bits_addr,
  input  [7:0]   io_req_bits_chosenWay,
  input          io_resp_ready,
  output         io_resp_valid,
  output [31:0]  io_resp_bits_data,
  output [31:0]  io_resp_bits_blockData_0,
  output [31:0]  io_resp_bits_blockData_1,
  output [31:0]  io_resp_bits_blockData_2,
  output [31:0]  io_resp_bits_blockData_3,
  output [31:0]  io_resp_bits_blockData_4,
  output [31:0]  io_resp_bits_blockData_5,
  output [31:0]  io_resp_bits_blockData_6,
  output [31:0]  io_resp_bits_blockData_7,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [31:0]  io_tlbus_req_bits_address,
  output         io_tlbus_resp_ready,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data,
  output         io_dirWrite_req_valid,
  output [31:0]  io_dirWrite_req_bits_addr,
  output [7:0]   io_dirWrite_req_bits_way,
  output         io_dataWrite_req_valid,
  output [6:0]   io_dataWrite_req_bits_set,
  output [31:0]  io_dataWrite_req_bits_data_0,
  output [31:0]  io_dataWrite_req_bits_data_1,
  output [31:0]  io_dataWrite_req_bits_data_2,
  output [31:0]  io_dataWrite_req_bits_data_3,
  output [31:0]  io_dataWrite_req_bits_data_4,
  output [31:0]  io_dataWrite_req_bits_data_5,
  output [31:0]  io_dataWrite_req_bits_data_6,
  output [31:0]  io_dataWrite_req_bits_data_7,
  output [7:0]   io_dataWrite_req_bits_blockMask,
  output [7:0]   io_dataWrite_req_bits_way
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[RefillPipe.scala 42:24]
  wire  _io_req_ready_T = state == 2'h0; // @[RefillPipe.scala 45:27]
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] reqReg_addr; // @[Reg.scala 19:16]
  reg [7:0] reqReg_chosenWay; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  reg  reqValidReg; // @[Reg.scala 19:16]
  wire  _GEN_2 = _reqReg_T | reqValidReg; // @[Reg.scala 19:16 20:{18,22}]
  wire [7:0] dataBlockSelOH = 8'h1 << reqReg_addr[4:2]; // @[OneHot.scala 57:35]
  reg  beatCounter_value; // @[Counter.scala 61:40]
  wire [1:0] beatOH = 2'h1 << beatCounter_value; // @[OneHot.scala 64:12]
  wire  _refillFire_T = io_tlbus_resp_ready & io_tlbus_resp_valid; // @[Decoupled.scala 51:35]
  wire  refillFire = _refillFire_T & io_tlbus_resp_bits_opcode == 3'h1; // @[RefillPipe.scala 59:41]
  wire  refillLastBeat = refillFire & beatCounter_value; // @[RefillPipe.scala 60:37]
  wire  _T_2 = io_tlbus_req_ready & io_tlbus_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_4 = _T_2 ? 2'h2 : {{1'd0}, _reqReg_T}; // @[RefillPipe.scala 71:33 72:23]
  wire  _GEN_5 = _T_2 ? 1'h0 : _GEN_2; // @[RefillPipe.scala 71:33 73:25]
  wire [1:0] _GEN_6 = _io_req_ready_T ? _GEN_4 : 2'h0; // @[RefillPipe.scala 66:27 43:29]
  wire  _GEN_7 = _io_req_ready_T ? _GEN_5 : _GEN_2; // @[RefillPipe.scala 66:27]
  wire [1:0] _GEN_8 = _T_2 ? 2'h2 : 2'h1; // @[RefillPipe.scala 80:19 81:33 82:23]
  wire  _T_5 = state == 2'h2; // @[RefillPipe.scala 89:16]
  wire  _T_6 = io_resp_ready & io_resp_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_12 = _T_6 ? 2'h0 : 2'h3; // @[RefillPipe.scala 92:23 93:32 94:27]
  wire  _T_7 = state == 2'h3; // @[RefillPipe.scala 105:16]
  wire  refillSafe = refillFire & _T_5; // @[RefillPipe.scala 115:33]
  wire [3:0] _blockMask_T_3 = beatOH[0] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _blockMask_T_5 = beatOH[1] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [255:0] _T_9 = {io_tlbus_resp_bits_data,io_tlbus_resp_bits_data}; // @[Cat.scala 33:92]
  reg [31:0] refillBlockDataArray_0_0; // @[RefillPipe.scala 133:39]
  reg [31:0] refillBlockDataArray_0_1; // @[RefillPipe.scala 133:39]
  reg [31:0] refillBlockDataArray_0_2; // @[RefillPipe.scala 133:39]
  reg [31:0] refillBlockDataArray_0_3; // @[RefillPipe.scala 133:39]
  wire [255:0] _io_resp_bits_data_T = {io_tlbus_resp_bits_data,refillBlockDataArray_0_3,refillBlockDataArray_0_2,
    refillBlockDataArray_0_1,refillBlockDataArray_0_0}; // @[RefillPipe.scala 141:72]
  wire [31:0] _io_resp_bits_data_T_17 = dataBlockSelOH[0] ? _io_resp_bits_data_T[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_18 = dataBlockSelOH[1] ? _io_resp_bits_data_T[63:32] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_19 = dataBlockSelOH[2] ? _io_resp_bits_data_T[95:64] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_20 = dataBlockSelOH[3] ? _io_resp_bits_data_T[127:96] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_21 = dataBlockSelOH[4] ? _io_resp_bits_data_T[159:128] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_22 = dataBlockSelOH[5] ? _io_resp_bits_data_T[191:160] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_23 = dataBlockSelOH[6] ? _io_resp_bits_data_T[223:192] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_24 = dataBlockSelOH[7] ? _io_resp_bits_data_T[255:224] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_25 = _io_resp_bits_data_T_17 | _io_resp_bits_data_T_18; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_26 = _io_resp_bits_data_T_25 | _io_resp_bits_data_T_19; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_27 = _io_resp_bits_data_T_26 | _io_resp_bits_data_T_20; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_28 = _io_resp_bits_data_T_27 | _io_resp_bits_data_T_21; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_29 = _io_resp_bits_data_T_28 | _io_resp_bits_data_T_22; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_30 = _io_resp_bits_data_T_29 | _io_resp_bits_data_T_23; // @[Mux.scala 27:73]
  assign io_req_ready = state == 2'h0; // @[RefillPipe.scala 45:27]
  assign io_resp_valid = _T_7 | refillLastBeat; // @[RefillPipe.scala 140:38]
  assign io_resp_bits_data = _io_resp_bits_data_T_30 | _io_resp_bits_data_T_24; // @[Mux.scala 27:73]
  assign io_resp_bits_blockData_0 = _io_resp_bits_data_T[31:0]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_1 = _io_resp_bits_data_T[63:32]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_2 = _io_resp_bits_data_T[95:64]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_3 = _io_resp_bits_data_T[127:96]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_4 = _io_resp_bits_data_T[159:128]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_5 = _io_resp_bits_data_T[191:160]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_6 = _io_resp_bits_data_T[223:192]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_7 = _io_resp_bits_data_T[255:224]; // @[RefillPipe.scala 142:55]
  assign io_tlbus_req_valid = _reqReg_T | reqValidReg; // @[RefillPipe.scala 50:23]
  assign io_tlbus_req_bits_address = {_GEN_0[31:5],5'h0}; // @[Cat.scala 33:92]
  assign io_tlbus_resp_ready = 1'h1; // @[RefillPipe.scala 62:51]
  assign io_dirWrite_req_valid = refillSafe & beatCounter_value; // @[RefillPipe.scala 116:41]
  assign io_dirWrite_req_bits_addr = reqReg_addr; // @[RefillPipe.scala 117:31]
  assign io_dirWrite_req_bits_way = reqReg_chosenWay; // @[RefillPipe.scala 122:30]
  assign io_dataWrite_req_valid = refillFire & _T_5; // @[RefillPipe.scala 115:33]
  assign io_dataWrite_req_bits_set = reqReg_addr[11:5]; // @[Parameters.scala 50:11]
  assign io_dataWrite_req_bits_data_0 = _T_9[31:0]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_1 = _T_9[63:32]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_2 = _T_9[95:64]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_3 = _T_9[127:96]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_4 = _T_9[159:128]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_5 = _T_9[191:160]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_6 = _T_9[223:192]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_7 = _T_9[255:224]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_blockMask = {_blockMask_T_5,_blockMask_T_3}; // @[Cat.scala 33:92]
  assign io_dataWrite_req_bits_way = reqReg_chosenWay; // @[RefillPipe.scala 128:31]
  always @(posedge clock) begin
    if (reset) begin // @[RefillPipe.scala 42:24]
      state <= 2'h0; // @[RefillPipe.scala 42:24]
    end else if (state == 2'h3) begin // @[RefillPipe.scala 105:27]
      state <= _GEN_12;
    end else if (state == 2'h2) begin // @[RefillPipe.scala 89:33]
      if (refillLastBeat) begin // @[RefillPipe.scala 91:30]
        state <= _GEN_12;
      end else begin
        state <= 2'h2;
      end
    end else if (state == 2'h1) begin // @[RefillPipe.scala 79:26]
      state <= _GEN_8;
    end else begin
      state <= _GEN_6;
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_addr <= io_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_chosenWay <= io_req_bits_chosenWay; // @[Reg.scala 20:22]
    end
    if (state == 2'h1) begin // @[RefillPipe.scala 79:26]
      if (_T_2) begin // @[RefillPipe.scala 81:33]
        reqValidReg <= 1'h0; // @[RefillPipe.scala 83:25]
      end else begin
        reqValidReg <= _GEN_7;
      end
    end else begin
      reqValidReg <= _GEN_7;
    end
    if (reset) begin // @[Counter.scala 61:40]
      beatCounter_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (state == 2'h2) begin // @[RefillPipe.scala 89:33]
      if (refillLastBeat) begin // @[RefillPipe.scala 91:30]
        beatCounter_value <= 1'h0; // @[Counter.scala 98:11]
      end else if (refillFire) begin // @[RefillPipe.scala 97:32]
        beatCounter_value <= beatCounter_value + 1'h1; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[RefillPipe.scala 133:39]
      refillBlockDataArray_0_0 <= 32'h0; // @[RefillPipe.scala 133:39]
    end else if (refillFire) begin // @[RefillPipe.scala 134:22]
      if (~beatCounter_value) begin // @[RefillPipe.scala 135:49]
        refillBlockDataArray_0_0 <= io_tlbus_resp_bits_data[31:0]; // @[RefillPipe.scala 135:49]
      end
    end
    if (reset) begin // @[RefillPipe.scala 133:39]
      refillBlockDataArray_0_1 <= 32'h0; // @[RefillPipe.scala 133:39]
    end else if (refillFire) begin // @[RefillPipe.scala 134:22]
      if (~beatCounter_value) begin // @[RefillPipe.scala 135:49]
        refillBlockDataArray_0_1 <= io_tlbus_resp_bits_data[63:32]; // @[RefillPipe.scala 135:49]
      end
    end
    if (reset) begin // @[RefillPipe.scala 133:39]
      refillBlockDataArray_0_2 <= 32'h0; // @[RefillPipe.scala 133:39]
    end else if (refillFire) begin // @[RefillPipe.scala 134:22]
      if (~beatCounter_value) begin // @[RefillPipe.scala 135:49]
        refillBlockDataArray_0_2 <= io_tlbus_resp_bits_data[95:64]; // @[RefillPipe.scala 135:49]
      end
    end
    if (reset) begin // @[RefillPipe.scala 133:39]
      refillBlockDataArray_0_3 <= 32'h0; // @[RefillPipe.scala 133:39]
    end else if (refillFire) begin // @[RefillPipe.scala 134:22]
      if (~beatCounter_value) begin // @[RefillPipe.scala 135:49]
        refillBlockDataArray_0_3 <= io_tlbus_resp_bits_data[127:96]; // @[RefillPipe.scala 135:49]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reqReg_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqReg_chosenWay = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  reqValidReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  beatCounter_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  refillBlockDataArray_0_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  refillBlockDataArray_0_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  refillBlockDataArray_0_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  refillBlockDataArray_0_3 = _RAND_8[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RefillBuffer(
  input          clock,
  input          reset,
  input          io_write_valid,
  input  [31:0]  io_write_bits_cacheLineAddr,
  input  [127:0] io_write_bits_data,
  output [31:0]  io_read_cacheLineAddr_0,
  output [31:0]  io_read_cacheLineAddr_1,
  output [31:0]  io_read_cacheLineData_0_0,
  output [31:0]  io_read_cacheLineData_0_1,
  output [31:0]  io_read_cacheLineData_0_2,
  output [31:0]  io_read_cacheLineData_0_3,
  output [31:0]  io_read_cacheLineData_0_4,
  output [31:0]  io_read_cacheLineData_0_5,
  output [31:0]  io_read_cacheLineData_0_6,
  output [31:0]  io_read_cacheLineData_0_7,
  output [31:0]  io_read_cacheLineData_1_0,
  output [31:0]  io_read_cacheLineData_1_1,
  output [31:0]  io_read_cacheLineData_1_2,
  output [31:0]  io_read_cacheLineData_1_3,
  output [31:0]  io_read_cacheLineData_1_4,
  output [31:0]  io_read_cacheLineData_1_5,
  output [31:0]  io_read_cacheLineData_1_6,
  output [31:0]  io_read_cacheLineData_1_7,
  output         io_read_valids_0,
  output         io_read_valids_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] buf_0_0; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_1; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_2; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_3; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_4; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_5; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_6; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_7; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_0; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_1; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_2; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_3; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_4; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_5; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_6; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_7; // @[RefillBuffer.scala 23:18]
  reg [31:0] addr_0; // @[RefillBuffer.scala 24:19]
  reg [31:0] addr_1; // @[RefillBuffer.scala 24:19]
  reg  wrPtr_value; // @[Counter.scala 61:40]
  reg  beatCounter_value; // @[Counter.scala 61:40]
  wire [31:0] _addr_T_2 = {io_write_bits_cacheLineAddr[31:5],5'h0}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_60 = {{1'd0}, beatCounter_value}; // @[RefillBuffer.scala 23:18 43:{45,45}]
  wire [2:0] _GEN_66 = {{2'd0}, beatCounter_value}; // @[RefillBuffer.scala 23:18 43:{45,45}]
  assign io_read_cacheLineAddr_0 = addr_0; // @[RefillBuffer.scala 47:27]
  assign io_read_cacheLineAddr_1 = addr_1; // @[RefillBuffer.scala 47:27]
  assign io_read_cacheLineData_0_0 = buf_0_0; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_1 = buf_0_1; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_2 = buf_0_2; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_3 = buf_0_3; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_4 = buf_0_4; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_5 = buf_0_5; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_6 = buf_0_6; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_7 = buf_0_7; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_0 = buf_1_0; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_1 = buf_1_1; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_2 = buf_1_2; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_3 = buf_1_3; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_4 = buf_1_4; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_5 = buf_1_5; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_6 = buf_1_6; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_7 = buf_1_7; // @[RefillBuffer.scala 48:27]
  assign io_read_valids_0 = 1'h0; // @[RefillBuffer.scala 49:20]
  assign io_read_valids_1 = 1'h0; // @[RefillBuffer.scala 49:20]
  always @(posedge clock) begin
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & ~beatCounter_value) begin // @[RefillBuffer.scala 43:45]
        buf_0_0 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & beatCounter_value) begin // @[RefillBuffer.scala 43:45]
        buf_0_1 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 2'h2 == _GEN_60) begin // @[RefillBuffer.scala 43:45]
        buf_0_2 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 2'h3 == _GEN_60) begin // @[RefillBuffer.scala 43:45]
        buf_0_3 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 3'h4 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_0_4 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 3'h5 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_0_5 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 3'h6 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_0_6 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 3'h7 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_0_7 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & ~beatCounter_value) begin // @[RefillBuffer.scala 43:45]
        buf_1_0 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & beatCounter_value) begin // @[RefillBuffer.scala 43:45]
        buf_1_1 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 2'h2 == _GEN_60) begin // @[RefillBuffer.scala 43:45]
        buf_1_2 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 2'h3 == _GEN_60) begin // @[RefillBuffer.scala 43:45]
        buf_1_3 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 3'h4 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_1_4 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 3'h5 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_1_5 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 3'h6 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_1_6 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 3'h7 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_1_7 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid & beatCounter_value) begin // @[RefillBuffer.scala 34:37]
      if (~wrPtr_value) begin // @[RefillBuffer.scala 37:27]
        addr_0 <= _addr_T_2; // @[RefillBuffer.scala 37:27]
      end
    end
    if (io_write_valid & beatCounter_value) begin // @[RefillBuffer.scala 34:37]
      if (wrPtr_value) begin // @[RefillBuffer.scala 37:27]
        addr_1 <= _addr_T_2; // @[RefillBuffer.scala 37:27]
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      wrPtr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (io_write_valid & beatCounter_value) begin // @[RefillBuffer.scala 34:37]
      wrPtr_value <= wrPtr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      beatCounter_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (io_write_valid & beatCounter_value) begin // @[RefillBuffer.scala 34:37]
      beatCounter_value <= 1'h0; // @[Counter.scala 98:11]
    end else if (io_write_valid) begin // @[RefillBuffer.scala 38:31]
      beatCounter_value <= beatCounter_value + 1'h1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buf_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  buf_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  buf_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  buf_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  buf_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  buf_0_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  buf_0_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  buf_0_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  buf_1_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  buf_1_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  buf_1_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  buf_1_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  buf_1_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  buf_1_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  buf_1_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  buf_1_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  addr_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  addr_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  wrPtr_value = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  beatCounter_value = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_data,
  input  [31:0] io_in_0_bits_addr,
  input  [31:0] io_in_0_bits_inst_0,
  input  [31:0] io_in_0_bits_inst_1,
  input  [31:0] io_in_0_bits_inst_2,
  input  [31:0] io_in_0_bits_inst_3,
  input  [2:0]  io_in_0_bits_size,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_data,
  input  [31:0] io_in_1_bits_addr,
  input  [31:0] io_in_1_bits_inst_0,
  input  [31:0] io_in_1_bits_inst_1,
  input  [31:0] io_in_1_bits_inst_2,
  input  [31:0] io_in_1_bits_inst_3,
  input  [2:0]  io_in_1_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_data,
  output [31:0] io_out_bits_addr,
  output [31:0] io_out_bits_inst_0,
  output [31:0] io_out_bits_inst_1,
  output [31:0] io_out_bits_inst_2,
  output [31:0] io_out_bits_inst_3,
  output [2:0]  io_out_bits_size
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_inst_0 = io_in_0_valid ? io_in_0_bits_inst_0 : io_in_1_bits_inst_0; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_inst_1 = io_in_0_valid ? io_in_0_bits_inst_1 : io_in_1_bits_inst_1; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_inst_2 = io_in_0_valid ? io_in_0_bits_inst_2 : io_in_1_bits_inst_2; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_inst_3 = io_in_0_valid ? io_in_0_bits_inst_3 : io_in_1_bits_inst_3; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_size = io_in_0_valid ? io_in_0_bits_size : io_in_1_bits_size; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module ICache(
  input          clock,
  input          reset,
  output         io_read_req_ready,
  input          io_read_req_valid,
  input  [31:0]  io_read_req_bits_addr,
  input          io_read_resp_ready,
  output         io_read_resp_valid,
  output [31:0]  io_read_resp_bits_data,
  output [31:0]  io_read_resp_bits_addr,
  output [31:0]  io_read_resp_bits_inst_0,
  output [31:0]  io_read_resp_bits_inst_1,
  output [31:0]  io_read_resp_bits_inst_2,
  output [31:0]  io_read_resp_bits_inst_3,
  output [2:0]   io_read_resp_bits_size,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [31:0]  io_tlbus_req_bits_address,
  output         io_tlbus_resp_ready,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
`endif // RANDOMIZE_REG_INIT
  wire  db_clock; // @[ICache.scala 59:20]
  wire  db_reset; // @[ICache.scala 59:20]
  wire  db_io_read_req_ready; // @[ICache.scala 59:20]
  wire  db_io_read_req_valid; // @[ICache.scala 59:20]
  wire [6:0] db_io_read_req_bits_set; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_0_0; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_0_1; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_0_2; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_0_3; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_0_4; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_0_5; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_0_6; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_0_7; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_1_0; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_1_1; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_1_2; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_1_3; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_1_4; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_1_5; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_1_6; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_1_7; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_2_0; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_2_1; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_2_2; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_2_3; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_2_4; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_2_5; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_2_6; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_2_7; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_3_0; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_3_1; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_3_2; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_3_3; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_3_4; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_3_5; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_3_6; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_3_7; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_4_0; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_4_1; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_4_2; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_4_3; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_4_4; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_4_5; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_4_6; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_4_7; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_5_0; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_5_1; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_5_2; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_5_3; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_5_4; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_5_5; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_5_6; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_5_7; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_6_0; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_6_1; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_6_2; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_6_3; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_6_4; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_6_5; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_6_6; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_6_7; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_7_0; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_7_1; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_7_2; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_7_3; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_7_4; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_7_5; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_7_6; // @[ICache.scala 59:20]
  wire [31:0] db_io_read_resp_7_7; // @[ICache.scala 59:20]
  wire  db_io_write_req_ready; // @[ICache.scala 59:20]
  wire  db_io_write_req_valid; // @[ICache.scala 59:20]
  wire [6:0] db_io_write_req_bits_set; // @[ICache.scala 59:20]
  wire [31:0] db_io_write_req_bits_data_0; // @[ICache.scala 59:20]
  wire [31:0] db_io_write_req_bits_data_1; // @[ICache.scala 59:20]
  wire [31:0] db_io_write_req_bits_data_2; // @[ICache.scala 59:20]
  wire [31:0] db_io_write_req_bits_data_3; // @[ICache.scala 59:20]
  wire [31:0] db_io_write_req_bits_data_4; // @[ICache.scala 59:20]
  wire [31:0] db_io_write_req_bits_data_5; // @[ICache.scala 59:20]
  wire [31:0] db_io_write_req_bits_data_6; // @[ICache.scala 59:20]
  wire [31:0] db_io_write_req_bits_data_7; // @[ICache.scala 59:20]
  wire [7:0] db_io_write_req_bits_blockMask; // @[ICache.scala 59:20]
  wire [7:0] db_io_write_req_bits_way; // @[ICache.scala 59:20]
  wire  dir_clock; // @[ICache.scala 60:21]
  wire  dir_reset; // @[ICache.scala 60:21]
  wire  dir_io_read_req_ready; // @[ICache.scala 60:21]
  wire  dir_io_read_req_valid; // @[ICache.scala 60:21]
  wire [31:0] dir_io_read_req_bits_addr; // @[ICache.scala 60:21]
  wire  dir_io_read_resp_bits_hit; // @[ICache.scala 60:21]
  wire [7:0] dir_io_read_resp_bits_chosenWay; // @[ICache.scala 60:21]
  wire  dir_io_write_req_ready; // @[ICache.scala 60:21]
  wire  dir_io_write_req_valid; // @[ICache.scala 60:21]
  wire [31:0] dir_io_write_req_bits_addr; // @[ICache.scala 60:21]
  wire [7:0] dir_io_write_req_bits_way; // @[ICache.scala 60:21]
  wire  refillPipe_clock; // @[ICache.scala 61:28]
  wire  refillPipe_reset; // @[ICache.scala 61:28]
  wire  refillPipe_io_req_ready; // @[ICache.scala 61:28]
  wire  refillPipe_io_req_valid; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_req_bits_addr; // @[ICache.scala 61:28]
  wire [7:0] refillPipe_io_req_bits_chosenWay; // @[ICache.scala 61:28]
  wire  refillPipe_io_resp_ready; // @[ICache.scala 61:28]
  wire  refillPipe_io_resp_valid; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_resp_bits_data; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_0; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_1; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_2; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_3; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_4; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_5; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_6; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_7; // @[ICache.scala 61:28]
  wire  refillPipe_io_tlbus_req_ready; // @[ICache.scala 61:28]
  wire  refillPipe_io_tlbus_req_valid; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_tlbus_req_bits_address; // @[ICache.scala 61:28]
  wire  refillPipe_io_tlbus_resp_ready; // @[ICache.scala 61:28]
  wire  refillPipe_io_tlbus_resp_valid; // @[ICache.scala 61:28]
  wire [2:0] refillPipe_io_tlbus_resp_bits_opcode; // @[ICache.scala 61:28]
  wire [127:0] refillPipe_io_tlbus_resp_bits_data; // @[ICache.scala 61:28]
  wire  refillPipe_io_dirWrite_req_valid; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_dirWrite_req_bits_addr; // @[ICache.scala 61:28]
  wire [7:0] refillPipe_io_dirWrite_req_bits_way; // @[ICache.scala 61:28]
  wire  refillPipe_io_dataWrite_req_valid; // @[ICache.scala 61:28]
  wire [6:0] refillPipe_io_dataWrite_req_bits_set; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_0; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_1; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_2; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_3; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_4; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_5; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_6; // @[ICache.scala 61:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_7; // @[ICache.scala 61:28]
  wire [7:0] refillPipe_io_dataWrite_req_bits_blockMask; // @[ICache.scala 61:28]
  wire [7:0] refillPipe_io_dataWrite_req_bits_way; // @[ICache.scala 61:28]
  wire  refillBuffer_clock; // @[ICache.scala 68:30]
  wire  refillBuffer_reset; // @[ICache.scala 68:30]
  wire  refillBuffer_io_write_valid; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_write_bits_cacheLineAddr; // @[ICache.scala 68:30]
  wire [127:0] refillBuffer_io_write_bits_data; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineAddr_0; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineAddr_1; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_0; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_1; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_2; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_3; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_4; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_5; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_6; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_7; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_0; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_1; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_2; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_3; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_4; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_5; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_6; // @[ICache.scala 68:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_7; // @[ICache.scala 68:30]
  wire  refillBuffer_io_read_valids_0; // @[ICache.scala 68:30]
  wire  refillBuffer_io_read_valids_1; // @[ICache.scala 68:30]
  wire  readRespArb_io_in_0_ready; // @[ICache.scala 212:29]
  wire  readRespArb_io_in_0_valid; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_0_bits_data; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_0_bits_addr; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_0_bits_inst_0; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_0_bits_inst_1; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_0_bits_inst_2; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_0_bits_inst_3; // @[ICache.scala 212:29]
  wire [2:0] readRespArb_io_in_0_bits_size; // @[ICache.scala 212:29]
  wire  readRespArb_io_in_1_ready; // @[ICache.scala 212:29]
  wire  readRespArb_io_in_1_valid; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_1_bits_data; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_1_bits_addr; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_1_bits_inst_0; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_1_bits_inst_1; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_1_bits_inst_2; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_in_1_bits_inst_3; // @[ICache.scala 212:29]
  wire [2:0] readRespArb_io_in_1_bits_size; // @[ICache.scala 212:29]
  wire  readRespArb_io_out_ready; // @[ICache.scala 212:29]
  wire  readRespArb_io_out_valid; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_out_bits_data; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_out_bits_addr; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_out_bits_inst_0; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_out_bits_inst_1; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_out_bits_inst_2; // @[ICache.scala 212:29]
  wire [31:0] readRespArb_io_out_bits_inst_3; // @[ICache.scala 212:29]
  wire [2:0] readRespArb_io_out_bits_size; // @[ICache.scala 212:29]
  reg  s0_full; // @[ICache.scala 78:26]
  wire  s0_latch = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  reg  s1_full; // @[ICache.scala 116:26]
  reg  s1_info_dirInfo_hit; // @[Reg.scala 19:16]
  wire  s1_resp_ready = readRespArb_io_in_1_ready; // @[ICache.scala 146:27 214:26]
  wire  _s1_resp_valid_T = ~s1_info_dirInfo_hit; // @[ICache.scala 147:47]
  reg [31:0] s1_info_req_addr; // @[Reg.scala 19:16]
  wire [31:0] _bypassVec_T_2 = {s1_info_req_addr[31:5],5'h0}; // @[Cat.scala 33:92]
  wire  bypassVec_0 = refillBuffer_io_read_cacheLineAddr_0 == _bypassVec_T_2 & refillBuffer_io_read_valids_0; // @[ICache.scala 128:154]
  wire  bypassVec_1 = refillBuffer_io_read_cacheLineAddr_1 == _bypassVec_T_2 & refillBuffer_io_read_valids_1; // @[ICache.scala 128:154]
  wire [1:0] _s1_bypass_T = {bypassVec_0,bypassVec_1}; // @[Cat.scala 33:92]
  wire  s1_bypass = |_s1_bypass_T & s1_full & _s1_resp_valid_T; // @[ICache.scala 129:51]
  wire  _s1_resp_valid_T_1 = ~s1_info_dirInfo_hit & s1_bypass; // @[ICache.scala 147:68]
  reg  s2_full; // @[ICache.scala 167:26]
  reg  s2_dirInfo_hit; // @[Reg.scala 19:16]
  reg  s2_bypass; // @[Reg.scala 19:16]
  wire  _s2_valid_T_1 = ~s2_dirInfo_hit; // @[ICache.scala 202:60]
  wire  s2_resp_ready = readRespArb_io_in_0_ready; // @[ICache.scala 192:27 213:26]
  wire  _s2_resp_valid_T_2 = refillPipe_io_resp_ready & refillPipe_io_resp_valid; // @[Decoupled.scala 51:35]
  reg  s2_refillValid; // @[ICache.scala 185:33]
  wire  _s2_resp_valid_T_3 = _s2_resp_valid_T_2 | s2_refillValid; // @[ICache.scala 193:77]
  wire  s2_resp_valid = _s2_valid_T_1 & s2_full & (_s2_resp_valid_T_2 | s2_refillValid); // @[ICache.scala 193:49]
  wire  _s2_valid_T_2 = s2_resp_ready & s2_resp_valid; // @[Decoupled.scala 51:35]
  wire  s2_fire = s2_full & (s2_dirInfo_hit | s2_bypass | ~s2_dirInfo_hit & _s2_valid_T_2); // @[ICache.scala 202:25]
  wire  s2_ready = ~s2_full | s2_fire; // @[ICache.scala 173:26]
  wire  s1_resp_valid = (s1_info_dirInfo_hit | ~s1_info_dirInfo_hit & s1_bypass) & s1_full & s2_ready; // @[ICache.scala 147:94]
  wire  _s1_valid_T = s1_resp_ready & s1_resp_valid; // @[Decoupled.scala 51:35]
  wire  _s1_valid_T_3 = refillPipe_io_req_ready & refillPipe_io_req_valid; // @[Decoupled.scala 51:35]
  wire  _s1_valid_T_5 = ~s1_bypass; // @[ICache.scala 156:75]
  wire  _s1_valid_T_6 = _s1_resp_valid_T & _s1_valid_T_3 & ~s1_bypass; // @[ICache.scala 156:72]
  wire  _s1_valid_T_7 = s1_info_dirInfo_hit & _s1_valid_T | _s1_valid_T_6; // @[ICache.scala 155:66]
  wire  _s1_valid_T_11 = _s1_resp_valid_T_1 & _s1_valid_T; // @[ICache.scala 157:59]
  wire  _s1_valid_T_12 = _s1_valid_T_7 | _s1_valid_T_11; // @[ICache.scala 156:86]
  wire  s1_valid = s1_full & _s1_valid_T_12; // @[ICache.scala 155:25]
  wire  s1_fire = s1_valid & s2_ready; // @[ICache.scala 118:28]
  wire  s1_ready = ~s1_full | s1_fire; // @[ICache.scala 123:26]
  wire  s0_fire = s0_full & s1_ready; // @[ICache.scala 80:28]
  reg [31:0] s0_req_r_addr; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = s0_latch ? io_read_req_bits_addr : s0_req_r_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_1 = s0_full & s0_fire ? 1'h0 : s0_full; // @[ICache.scala 78:26 86:{35,45}]
  wire  _GEN_2 = s0_latch | _GEN_1; // @[ICache.scala 85:{20,30}]
  reg [7:0] s1_info_dirInfo_chosenWay; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_7; // @[Reg.scala 19:16]
  wire [31:0] s0_info_rdData_0_0 = db_io_read_resp_0_0; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_0_1 = db_io_read_resp_0_1; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_0_2 = db_io_read_resp_0_2; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_0_3 = db_io_read_resp_0_3; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_0_4 = db_io_read_resp_0_4; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_0_5 = db_io_read_resp_0_5; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_0_6 = db_io_read_resp_0_6; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_0_7 = db_io_read_resp_0_7; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_1_0 = db_io_read_resp_1_0; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_1_1 = db_io_read_resp_1_1; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_1_2 = db_io_read_resp_1_2; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_1_3 = db_io_read_resp_1_3; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_1_4 = db_io_read_resp_1_4; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_1_5 = db_io_read_resp_1_5; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_1_6 = db_io_read_resp_1_6; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_1_7 = db_io_read_resp_1_7; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_2_0 = db_io_read_resp_2_0; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_2_1 = db_io_read_resp_2_1; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_2_2 = db_io_read_resp_2_2; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_2_3 = db_io_read_resp_2_3; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_2_4 = db_io_read_resp_2_4; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_2_5 = db_io_read_resp_2_5; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_2_6 = db_io_read_resp_2_6; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_2_7 = db_io_read_resp_2_7; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_3_0 = db_io_read_resp_3_0; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_3_1 = db_io_read_resp_3_1; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_3_2 = db_io_read_resp_3_2; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_3_3 = db_io_read_resp_3_3; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_3_4 = db_io_read_resp_3_4; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_3_5 = db_io_read_resp_3_5; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_3_6 = db_io_read_resp_3_6; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_3_7 = db_io_read_resp_3_7; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_4_0 = db_io_read_resp_4_0; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_4_1 = db_io_read_resp_4_1; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_4_2 = db_io_read_resp_4_2; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_4_3 = db_io_read_resp_4_3; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_4_4 = db_io_read_resp_4_4; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_4_5 = db_io_read_resp_4_5; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_4_6 = db_io_read_resp_4_6; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_4_7 = db_io_read_resp_4_7; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_5_0 = db_io_read_resp_5_0; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_5_1 = db_io_read_resp_5_1; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_5_2 = db_io_read_resp_5_2; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_5_3 = db_io_read_resp_5_3; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_5_4 = db_io_read_resp_5_4; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_5_5 = db_io_read_resp_5_5; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_5_6 = db_io_read_resp_5_6; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_5_7 = db_io_read_resp_5_7; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_6_0 = db_io_read_resp_6_0; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_6_1 = db_io_read_resp_6_1; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_6_2 = db_io_read_resp_6_2; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_6_3 = db_io_read_resp_6_3; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_6_4 = db_io_read_resp_6_4; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_6_5 = db_io_read_resp_6_5; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_6_6 = db_io_read_resp_6_6; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_6_7 = db_io_read_resp_6_7; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_7_0 = db_io_read_resp_7_0; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_7_1 = db_io_read_resp_7_1; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_7_2 = db_io_read_resp_7_2; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_7_3 = db_io_read_resp_7_3; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_7_4 = db_io_read_resp_7_4; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_7_5 = db_io_read_resp_7_5; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_7_6 = db_io_read_resp_7_6; // @[ICache.scala 107:23 110:20]
  wire [31:0] s0_info_rdData_7_7 = db_io_read_resp_7_7; // @[ICache.scala 107:23 110:20]
  wire  s0_info_dirInfo_hit = dir_io_read_resp_bits_hit; // @[ICache.scala 107:23 108:21]
  wire [7:0] s0_info_dirInfo_chosenWay = dir_io_read_resp_bits_chosenWay; // @[ICache.scala 107:23 108:21]
  wire [7:0] s1_blockSel = 8'h1 << s1_info_req_addr[4:2]; // @[OneHot.scala 57:35]
  wire [31:0] _s1_rdBlockData_T_8 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_9 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_10 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_11 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_12 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_13 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_14 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_15 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_16 = _s1_rdBlockData_T_8 | _s1_rdBlockData_T_9; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_17 = _s1_rdBlockData_T_16 | _s1_rdBlockData_T_10; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_18 = _s1_rdBlockData_T_17 | _s1_rdBlockData_T_11; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_19 = _s1_rdBlockData_T_18 | _s1_rdBlockData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_20 = _s1_rdBlockData_T_19 | _s1_rdBlockData_T_13; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_21 = _s1_rdBlockData_T_20 | _s1_rdBlockData_T_14; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_0 = _s1_rdBlockData_T_21 | _s1_rdBlockData_T_15; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_23 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_24 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_25 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_26 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_27 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_28 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_29 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_30 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_31 = _s1_rdBlockData_T_23 | _s1_rdBlockData_T_24; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_32 = _s1_rdBlockData_T_31 | _s1_rdBlockData_T_25; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_33 = _s1_rdBlockData_T_32 | _s1_rdBlockData_T_26; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_34 = _s1_rdBlockData_T_33 | _s1_rdBlockData_T_27; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_35 = _s1_rdBlockData_T_34 | _s1_rdBlockData_T_28; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_36 = _s1_rdBlockData_T_35 | _s1_rdBlockData_T_29; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_1 = _s1_rdBlockData_T_36 | _s1_rdBlockData_T_30; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_38 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_39 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_40 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_41 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_42 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_43 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_44 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_45 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_46 = _s1_rdBlockData_T_38 | _s1_rdBlockData_T_39; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_47 = _s1_rdBlockData_T_46 | _s1_rdBlockData_T_40; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_48 = _s1_rdBlockData_T_47 | _s1_rdBlockData_T_41; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_49 = _s1_rdBlockData_T_48 | _s1_rdBlockData_T_42; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_50 = _s1_rdBlockData_T_49 | _s1_rdBlockData_T_43; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_51 = _s1_rdBlockData_T_50 | _s1_rdBlockData_T_44; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_2 = _s1_rdBlockData_T_51 | _s1_rdBlockData_T_45; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_53 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_54 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_55 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_56 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_57 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_58 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_59 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_60 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_61 = _s1_rdBlockData_T_53 | _s1_rdBlockData_T_54; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_62 = _s1_rdBlockData_T_61 | _s1_rdBlockData_T_55; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_63 = _s1_rdBlockData_T_62 | _s1_rdBlockData_T_56; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_64 = _s1_rdBlockData_T_63 | _s1_rdBlockData_T_57; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_65 = _s1_rdBlockData_T_64 | _s1_rdBlockData_T_58; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_66 = _s1_rdBlockData_T_65 | _s1_rdBlockData_T_59; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_3 = _s1_rdBlockData_T_66 | _s1_rdBlockData_T_60; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_68 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_69 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_70 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_71 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_72 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_73 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_74 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_75 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_76 = _s1_rdBlockData_T_68 | _s1_rdBlockData_T_69; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_77 = _s1_rdBlockData_T_76 | _s1_rdBlockData_T_70; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_78 = _s1_rdBlockData_T_77 | _s1_rdBlockData_T_71; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_79 = _s1_rdBlockData_T_78 | _s1_rdBlockData_T_72; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_80 = _s1_rdBlockData_T_79 | _s1_rdBlockData_T_73; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_81 = _s1_rdBlockData_T_80 | _s1_rdBlockData_T_74; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_4 = _s1_rdBlockData_T_81 | _s1_rdBlockData_T_75; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_83 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_84 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_85 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_86 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_87 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_88 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_89 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_90 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_91 = _s1_rdBlockData_T_83 | _s1_rdBlockData_T_84; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_92 = _s1_rdBlockData_T_91 | _s1_rdBlockData_T_85; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_93 = _s1_rdBlockData_T_92 | _s1_rdBlockData_T_86; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_94 = _s1_rdBlockData_T_93 | _s1_rdBlockData_T_87; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_95 = _s1_rdBlockData_T_94 | _s1_rdBlockData_T_88; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_96 = _s1_rdBlockData_T_95 | _s1_rdBlockData_T_89; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_5 = _s1_rdBlockData_T_96 | _s1_rdBlockData_T_90; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_98 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_99 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_100 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_101 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_102 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_103 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_104 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_105 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_106 = _s1_rdBlockData_T_98 | _s1_rdBlockData_T_99; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_107 = _s1_rdBlockData_T_106 | _s1_rdBlockData_T_100; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_108 = _s1_rdBlockData_T_107 | _s1_rdBlockData_T_101; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_109 = _s1_rdBlockData_T_108 | _s1_rdBlockData_T_102; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_110 = _s1_rdBlockData_T_109 | _s1_rdBlockData_T_103; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_111 = _s1_rdBlockData_T_110 | _s1_rdBlockData_T_104; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_6 = _s1_rdBlockData_T_111 | _s1_rdBlockData_T_105; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_113 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_114 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_115 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_116 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_117 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_118 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_119 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_120 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_121 = _s1_rdBlockData_T_113 | _s1_rdBlockData_T_114; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_122 = _s1_rdBlockData_T_121 | _s1_rdBlockData_T_115; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_123 = _s1_rdBlockData_T_122 | _s1_rdBlockData_T_116; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_124 = _s1_rdBlockData_T_123 | _s1_rdBlockData_T_117; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_125 = _s1_rdBlockData_T_124 | _s1_rdBlockData_T_118; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_126 = _s1_rdBlockData_T_125 | _s1_rdBlockData_T_119; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_7 = _s1_rdBlockData_T_126 | _s1_rdBlockData_T_120; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_8 = s1_blockSel[0] ? s1_rdBlockData_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_9 = s1_blockSel[1] ? s1_rdBlockData_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_10 = s1_blockSel[2] ? s1_rdBlockData_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_11 = s1_blockSel[3] ? s1_rdBlockData_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_12 = s1_blockSel[4] ? s1_rdBlockData_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_13 = s1_blockSel[5] ? s1_rdBlockData_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_14 = s1_blockSel[6] ? s1_rdBlockData_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_15 = s1_blockSel[7] ? s1_rdBlockData_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_16 = _s1_rdHitData_T_8 | _s1_rdHitData_T_9; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_17 = _s1_rdHitData_T_16 | _s1_rdHitData_T_10; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_18 = _s1_rdHitData_T_17 | _s1_rdHitData_T_11; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_19 = _s1_rdHitData_T_18 | _s1_rdHitData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_20 = _s1_rdHitData_T_19 | _s1_rdHitData_T_13; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_21 = _s1_rdHitData_T_20 | _s1_rdHitData_T_14; // @[Mux.scala 27:73]
  wire [31:0] s1_rdHitData = _s1_rdHitData_T_21 | _s1_rdHitData_T_15; // @[Mux.scala 27:73]
  wire  _GEN_79 = s1_full & s1_fire ? 1'h0 : s1_full; // @[ICache.scala 116:26 126:{35,45}]
  wire  _GEN_80 = s0_fire | _GEN_79; // @[ICache.scala 125:{20,30}]
  wire [1:0] _s1_bypassIdx_T = {bypassVec_1,bypassVec_0}; // @[Cat.scala 33:92]
  wire  s1_bypassIdx = _s1_bypassIdx_T[1]; // @[CircuitMath.scala 28:8]
  wire [31:0] _GEN_81 = refillBuffer_io_read_cacheLineData_0_0; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_82 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_0 : _GEN_81; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_8 = s1_blockSel[0] ? _GEN_82 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_83 = refillBuffer_io_read_cacheLineData_0_1; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_84 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_1 : _GEN_83; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_9 = s1_blockSel[1] ? _GEN_84 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_85 = refillBuffer_io_read_cacheLineData_0_2; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_86 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_2 : _GEN_85; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_10 = s1_blockSel[2] ? _GEN_86 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_87 = refillBuffer_io_read_cacheLineData_0_3; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_88 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_3 : _GEN_87; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_11 = s1_blockSel[3] ? _GEN_88 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_89 = refillBuffer_io_read_cacheLineData_0_4; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_90 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_4 : _GEN_89; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_12 = s1_blockSel[4] ? _GEN_90 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_91 = refillBuffer_io_read_cacheLineData_0_5; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_92 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_5 : _GEN_91; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_13 = s1_blockSel[5] ? _GEN_92 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_93 = refillBuffer_io_read_cacheLineData_0_6; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_94 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_6 : _GEN_93; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_14 = s1_blockSel[6] ? _GEN_94 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_95 = refillBuffer_io_read_cacheLineData_0_7; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_96 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_7 : _GEN_95; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_15 = s1_blockSel[7] ? _GEN_96 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_16 = _s1_bypassData_T_8 | _s1_bypassData_T_9; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_17 = _s1_bypassData_T_16 | _s1_bypassData_T_10; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_18 = _s1_bypassData_T_17 | _s1_bypassData_T_11; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_19 = _s1_bypassData_T_18 | _s1_bypassData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_20 = _s1_bypassData_T_19 | _s1_bypassData_T_13; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_21 = _s1_bypassData_T_20 | _s1_bypassData_T_14; // @[Mux.scala 27:73]
  wire [3:0] rdThreshole = 4'h8 - 4'h4; // @[ICache.scala 140:41]
  wire [2:0] s1_off = s1_info_req_addr[4:2]; // @[ICache.scala 141:34]
  wire [3:0] _GEN_116 = {{1'd0}, s1_info_req_addr[4:2]}; // @[ICache.scala 143:37]
  wire [3:0] _s1_respHitSize_T_2 = 4'h8 - _GEN_116; // @[ICache.scala 143:71]
  wire [3:0] s1_respHitSize = _GEN_116 >= rdThreshole ? _s1_respHitSize_T_2 : 4'h4; // @[ICache.scala 143:29]
  wire [255:0] _s1_respHitInst_T = {s1_rdBlockData_7,s1_rdBlockData_6,s1_rdBlockData_5,s1_rdBlockData_4,s1_rdBlockData_3
    ,s1_rdBlockData_2,s1_rdBlockData_1,s1_rdBlockData_0}; // @[ICache.scala 144:42]
  wire [7:0] _s1_respHitInst_T_1 = {s1_info_req_addr[4:2], 5'h0}; // @[ICache.scala 144:60]
  wire [255:0] _s1_respHitInst_T_2 = _s1_respHitInst_T >> _s1_respHitInst_T_1; // @[ICache.scala 144:49]
  wire [31:0] s1_respHitInst_0 = _s1_respHitInst_T_2[31:0]; // @[ICache.scala 144:111]
  wire [31:0] s1_respHitInst_1 = _s1_respHitInst_T_2[63:32]; // @[ICache.scala 144:111]
  wire [31:0] s1_respHitInst_2 = _s1_respHitInst_T_2[95:64]; // @[ICache.scala 144:111]
  wire [31:0] s1_respHitInst_3 = _s1_respHitInst_T_2[127:96]; // @[ICache.scala 144:111]
  wire [255:0] _s1_respBypassInst_T = {_GEN_96,_GEN_94,_GEN_92,_GEN_90,_GEN_88,_GEN_86,_GEN_84,_GEN_82}; // @[ICache.scala 145:49]
  wire [255:0] _s1_respBypassInst_T_2 = _s1_respBypassInst_T >> _s1_respHitInst_T_1; // @[ICache.scala 145:56]
  wire [31:0] s1_respBypassInst_0 = _s1_respBypassInst_T_2[31:0]; // @[ICache.scala 145:118]
  wire [31:0] s1_respBypassInst_1 = _s1_respBypassInst_T_2[63:32]; // @[ICache.scala 145:118]
  wire [31:0] s1_respBypassInst_2 = _s1_respBypassInst_T_2[95:64]; // @[ICache.scala 145:118]
  wire [31:0] s1_respBypassInst_3 = _s1_respBypassInst_T_2[127:96]; // @[ICache.scala 145:118]
  wire [31:0] s1_bypassData = _s1_bypassData_T_21 | _s1_bypassData_T_15; // @[Mux.scala 27:73]
  reg [31:0] s2_addr; // @[Reg.scala 19:16]
  wire  _GEN_110 = s2_full & s2_fire ? 1'h0 : s2_full; // @[ICache.scala 167:26 176:{35,45}]
  wire  _GEN_111 = s1_fire | _GEN_110; // @[ICache.scala 175:{20,30}]
  wire  _refillBuffer_io_write_valid_T = io_tlbus_resp_ready & io_tlbus_resp_valid; // @[Decoupled.scala 51:35]
  wire [2:0] s2_off = s2_addr[4:2]; // @[ICache.scala 189:25]
  wire [3:0] _GEN_118 = {{1'd0}, s2_off}; // @[ICache.scala 190:38]
  wire [3:0] _s2_respMissSize_T_2 = 4'h8 - _GEN_118; // @[ICache.scala 190:72]
  wire [3:0] s2_respMissSize = _GEN_118 >= rdThreshole ? _s2_respMissSize_T_2 : 4'h4; // @[ICache.scala 190:30]
  wire [255:0] _s2_respRefillInst_T = {refillPipe_io_resp_bits_blockData_7,refillPipe_io_resp_bits_blockData_6,
    refillPipe_io_resp_bits_blockData_5,refillPipe_io_resp_bits_blockData_4,refillPipe_io_resp_bits_blockData_3,
    refillPipe_io_resp_bits_blockData_2,refillPipe_io_resp_bits_blockData_1,refillPipe_io_resp_bits_blockData_0}; // @[ICache.scala 191:64]
  wire [7:0] _s2_respRefillInst_T_1 = {s2_off, 5'h0}; // @[ICache.scala 191:82]
  wire [255:0] _s2_respRefillInst_T_2 = _s2_respRefillInst_T >> _s2_respRefillInst_T_1; // @[ICache.scala 191:71]
  DataBankArray db ( // @[ICache.scala 59:20]
    .clock(db_clock),
    .reset(db_reset),
    .io_read_req_ready(db_io_read_req_ready),
    .io_read_req_valid(db_io_read_req_valid),
    .io_read_req_bits_set(db_io_read_req_bits_set),
    .io_read_resp_0_0(db_io_read_resp_0_0),
    .io_read_resp_0_1(db_io_read_resp_0_1),
    .io_read_resp_0_2(db_io_read_resp_0_2),
    .io_read_resp_0_3(db_io_read_resp_0_3),
    .io_read_resp_0_4(db_io_read_resp_0_4),
    .io_read_resp_0_5(db_io_read_resp_0_5),
    .io_read_resp_0_6(db_io_read_resp_0_6),
    .io_read_resp_0_7(db_io_read_resp_0_7),
    .io_read_resp_1_0(db_io_read_resp_1_0),
    .io_read_resp_1_1(db_io_read_resp_1_1),
    .io_read_resp_1_2(db_io_read_resp_1_2),
    .io_read_resp_1_3(db_io_read_resp_1_3),
    .io_read_resp_1_4(db_io_read_resp_1_4),
    .io_read_resp_1_5(db_io_read_resp_1_5),
    .io_read_resp_1_6(db_io_read_resp_1_6),
    .io_read_resp_1_7(db_io_read_resp_1_7),
    .io_read_resp_2_0(db_io_read_resp_2_0),
    .io_read_resp_2_1(db_io_read_resp_2_1),
    .io_read_resp_2_2(db_io_read_resp_2_2),
    .io_read_resp_2_3(db_io_read_resp_2_3),
    .io_read_resp_2_4(db_io_read_resp_2_4),
    .io_read_resp_2_5(db_io_read_resp_2_5),
    .io_read_resp_2_6(db_io_read_resp_2_6),
    .io_read_resp_2_7(db_io_read_resp_2_7),
    .io_read_resp_3_0(db_io_read_resp_3_0),
    .io_read_resp_3_1(db_io_read_resp_3_1),
    .io_read_resp_3_2(db_io_read_resp_3_2),
    .io_read_resp_3_3(db_io_read_resp_3_3),
    .io_read_resp_3_4(db_io_read_resp_3_4),
    .io_read_resp_3_5(db_io_read_resp_3_5),
    .io_read_resp_3_6(db_io_read_resp_3_6),
    .io_read_resp_3_7(db_io_read_resp_3_7),
    .io_read_resp_4_0(db_io_read_resp_4_0),
    .io_read_resp_4_1(db_io_read_resp_4_1),
    .io_read_resp_4_2(db_io_read_resp_4_2),
    .io_read_resp_4_3(db_io_read_resp_4_3),
    .io_read_resp_4_4(db_io_read_resp_4_4),
    .io_read_resp_4_5(db_io_read_resp_4_5),
    .io_read_resp_4_6(db_io_read_resp_4_6),
    .io_read_resp_4_7(db_io_read_resp_4_7),
    .io_read_resp_5_0(db_io_read_resp_5_0),
    .io_read_resp_5_1(db_io_read_resp_5_1),
    .io_read_resp_5_2(db_io_read_resp_5_2),
    .io_read_resp_5_3(db_io_read_resp_5_3),
    .io_read_resp_5_4(db_io_read_resp_5_4),
    .io_read_resp_5_5(db_io_read_resp_5_5),
    .io_read_resp_5_6(db_io_read_resp_5_6),
    .io_read_resp_5_7(db_io_read_resp_5_7),
    .io_read_resp_6_0(db_io_read_resp_6_0),
    .io_read_resp_6_1(db_io_read_resp_6_1),
    .io_read_resp_6_2(db_io_read_resp_6_2),
    .io_read_resp_6_3(db_io_read_resp_6_3),
    .io_read_resp_6_4(db_io_read_resp_6_4),
    .io_read_resp_6_5(db_io_read_resp_6_5),
    .io_read_resp_6_6(db_io_read_resp_6_6),
    .io_read_resp_6_7(db_io_read_resp_6_7),
    .io_read_resp_7_0(db_io_read_resp_7_0),
    .io_read_resp_7_1(db_io_read_resp_7_1),
    .io_read_resp_7_2(db_io_read_resp_7_2),
    .io_read_resp_7_3(db_io_read_resp_7_3),
    .io_read_resp_7_4(db_io_read_resp_7_4),
    .io_read_resp_7_5(db_io_read_resp_7_5),
    .io_read_resp_7_6(db_io_read_resp_7_6),
    .io_read_resp_7_7(db_io_read_resp_7_7),
    .io_write_req_ready(db_io_write_req_ready),
    .io_write_req_valid(db_io_write_req_valid),
    .io_write_req_bits_set(db_io_write_req_bits_set),
    .io_write_req_bits_data_0(db_io_write_req_bits_data_0),
    .io_write_req_bits_data_1(db_io_write_req_bits_data_1),
    .io_write_req_bits_data_2(db_io_write_req_bits_data_2),
    .io_write_req_bits_data_3(db_io_write_req_bits_data_3),
    .io_write_req_bits_data_4(db_io_write_req_bits_data_4),
    .io_write_req_bits_data_5(db_io_write_req_bits_data_5),
    .io_write_req_bits_data_6(db_io_write_req_bits_data_6),
    .io_write_req_bits_data_7(db_io_write_req_bits_data_7),
    .io_write_req_bits_blockMask(db_io_write_req_bits_blockMask),
    .io_write_req_bits_way(db_io_write_req_bits_way)
  );
  DCacheDirectory dir ( // @[ICache.scala 60:21]
    .clock(dir_clock),
    .reset(dir_reset),
    .io_read_req_ready(dir_io_read_req_ready),
    .io_read_req_valid(dir_io_read_req_valid),
    .io_read_req_bits_addr(dir_io_read_req_bits_addr),
    .io_read_resp_bits_hit(dir_io_read_resp_bits_hit),
    .io_read_resp_bits_chosenWay(dir_io_read_resp_bits_chosenWay),
    .io_write_req_ready(dir_io_write_req_ready),
    .io_write_req_valid(dir_io_write_req_valid),
    .io_write_req_bits_addr(dir_io_write_req_bits_addr),
    .io_write_req_bits_way(dir_io_write_req_bits_way)
  );
  RefillPipe refillPipe ( // @[ICache.scala 61:28]
    .clock(refillPipe_clock),
    .reset(refillPipe_reset),
    .io_req_ready(refillPipe_io_req_ready),
    .io_req_valid(refillPipe_io_req_valid),
    .io_req_bits_addr(refillPipe_io_req_bits_addr),
    .io_req_bits_chosenWay(refillPipe_io_req_bits_chosenWay),
    .io_resp_ready(refillPipe_io_resp_ready),
    .io_resp_valid(refillPipe_io_resp_valid),
    .io_resp_bits_data(refillPipe_io_resp_bits_data),
    .io_resp_bits_blockData_0(refillPipe_io_resp_bits_blockData_0),
    .io_resp_bits_blockData_1(refillPipe_io_resp_bits_blockData_1),
    .io_resp_bits_blockData_2(refillPipe_io_resp_bits_blockData_2),
    .io_resp_bits_blockData_3(refillPipe_io_resp_bits_blockData_3),
    .io_resp_bits_blockData_4(refillPipe_io_resp_bits_blockData_4),
    .io_resp_bits_blockData_5(refillPipe_io_resp_bits_blockData_5),
    .io_resp_bits_blockData_6(refillPipe_io_resp_bits_blockData_6),
    .io_resp_bits_blockData_7(refillPipe_io_resp_bits_blockData_7),
    .io_tlbus_req_ready(refillPipe_io_tlbus_req_ready),
    .io_tlbus_req_valid(refillPipe_io_tlbus_req_valid),
    .io_tlbus_req_bits_address(refillPipe_io_tlbus_req_bits_address),
    .io_tlbus_resp_ready(refillPipe_io_tlbus_resp_ready),
    .io_tlbus_resp_valid(refillPipe_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(refillPipe_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(refillPipe_io_tlbus_resp_bits_data),
    .io_dirWrite_req_valid(refillPipe_io_dirWrite_req_valid),
    .io_dirWrite_req_bits_addr(refillPipe_io_dirWrite_req_bits_addr),
    .io_dirWrite_req_bits_way(refillPipe_io_dirWrite_req_bits_way),
    .io_dataWrite_req_valid(refillPipe_io_dataWrite_req_valid),
    .io_dataWrite_req_bits_set(refillPipe_io_dataWrite_req_bits_set),
    .io_dataWrite_req_bits_data_0(refillPipe_io_dataWrite_req_bits_data_0),
    .io_dataWrite_req_bits_data_1(refillPipe_io_dataWrite_req_bits_data_1),
    .io_dataWrite_req_bits_data_2(refillPipe_io_dataWrite_req_bits_data_2),
    .io_dataWrite_req_bits_data_3(refillPipe_io_dataWrite_req_bits_data_3),
    .io_dataWrite_req_bits_data_4(refillPipe_io_dataWrite_req_bits_data_4),
    .io_dataWrite_req_bits_data_5(refillPipe_io_dataWrite_req_bits_data_5),
    .io_dataWrite_req_bits_data_6(refillPipe_io_dataWrite_req_bits_data_6),
    .io_dataWrite_req_bits_data_7(refillPipe_io_dataWrite_req_bits_data_7),
    .io_dataWrite_req_bits_blockMask(refillPipe_io_dataWrite_req_bits_blockMask),
    .io_dataWrite_req_bits_way(refillPipe_io_dataWrite_req_bits_way)
  );
  RefillBuffer refillBuffer ( // @[ICache.scala 68:30]
    .clock(refillBuffer_clock),
    .reset(refillBuffer_reset),
    .io_write_valid(refillBuffer_io_write_valid),
    .io_write_bits_cacheLineAddr(refillBuffer_io_write_bits_cacheLineAddr),
    .io_write_bits_data(refillBuffer_io_write_bits_data),
    .io_read_cacheLineAddr_0(refillBuffer_io_read_cacheLineAddr_0),
    .io_read_cacheLineAddr_1(refillBuffer_io_read_cacheLineAddr_1),
    .io_read_cacheLineData_0_0(refillBuffer_io_read_cacheLineData_0_0),
    .io_read_cacheLineData_0_1(refillBuffer_io_read_cacheLineData_0_1),
    .io_read_cacheLineData_0_2(refillBuffer_io_read_cacheLineData_0_2),
    .io_read_cacheLineData_0_3(refillBuffer_io_read_cacheLineData_0_3),
    .io_read_cacheLineData_0_4(refillBuffer_io_read_cacheLineData_0_4),
    .io_read_cacheLineData_0_5(refillBuffer_io_read_cacheLineData_0_5),
    .io_read_cacheLineData_0_6(refillBuffer_io_read_cacheLineData_0_6),
    .io_read_cacheLineData_0_7(refillBuffer_io_read_cacheLineData_0_7),
    .io_read_cacheLineData_1_0(refillBuffer_io_read_cacheLineData_1_0),
    .io_read_cacheLineData_1_1(refillBuffer_io_read_cacheLineData_1_1),
    .io_read_cacheLineData_1_2(refillBuffer_io_read_cacheLineData_1_2),
    .io_read_cacheLineData_1_3(refillBuffer_io_read_cacheLineData_1_3),
    .io_read_cacheLineData_1_4(refillBuffer_io_read_cacheLineData_1_4),
    .io_read_cacheLineData_1_5(refillBuffer_io_read_cacheLineData_1_5),
    .io_read_cacheLineData_1_6(refillBuffer_io_read_cacheLineData_1_6),
    .io_read_cacheLineData_1_7(refillBuffer_io_read_cacheLineData_1_7),
    .io_read_valids_0(refillBuffer_io_read_valids_0),
    .io_read_valids_1(refillBuffer_io_read_valids_1)
  );
  Arbiter readRespArb ( // @[ICache.scala 212:29]
    .io_in_0_ready(readRespArb_io_in_0_ready),
    .io_in_0_valid(readRespArb_io_in_0_valid),
    .io_in_0_bits_data(readRespArb_io_in_0_bits_data),
    .io_in_0_bits_addr(readRespArb_io_in_0_bits_addr),
    .io_in_0_bits_inst_0(readRespArb_io_in_0_bits_inst_0),
    .io_in_0_bits_inst_1(readRespArb_io_in_0_bits_inst_1),
    .io_in_0_bits_inst_2(readRespArb_io_in_0_bits_inst_2),
    .io_in_0_bits_inst_3(readRespArb_io_in_0_bits_inst_3),
    .io_in_0_bits_size(readRespArb_io_in_0_bits_size),
    .io_in_1_ready(readRespArb_io_in_1_ready),
    .io_in_1_valid(readRespArb_io_in_1_valid),
    .io_in_1_bits_data(readRespArb_io_in_1_bits_data),
    .io_in_1_bits_addr(readRespArb_io_in_1_bits_addr),
    .io_in_1_bits_inst_0(readRespArb_io_in_1_bits_inst_0),
    .io_in_1_bits_inst_1(readRespArb_io_in_1_bits_inst_1),
    .io_in_1_bits_inst_2(readRespArb_io_in_1_bits_inst_2),
    .io_in_1_bits_inst_3(readRespArb_io_in_1_bits_inst_3),
    .io_in_1_bits_size(readRespArb_io_in_1_bits_size),
    .io_out_ready(readRespArb_io_out_ready),
    .io_out_valid(readRespArb_io_out_valid),
    .io_out_bits_data(readRespArb_io_out_bits_data),
    .io_out_bits_addr(readRespArb_io_out_bits_addr),
    .io_out_bits_inst_0(readRespArb_io_out_bits_inst_0),
    .io_out_bits_inst_1(readRespArb_io_out_bits_inst_1),
    .io_out_bits_inst_2(readRespArb_io_out_bits_inst_2),
    .io_out_bits_inst_3(readRespArb_io_out_bits_inst_3),
    .io_out_bits_size(readRespArb_io_out_bits_size)
  );
  assign io_read_req_ready = ~s0_full; // @[ICache.scala 83:26]
  assign io_read_resp_valid = readRespArb_io_out_valid; // @[ICache.scala 215:18]
  assign io_read_resp_bits_data = readRespArb_io_out_bits_data; // @[ICache.scala 215:18]
  assign io_read_resp_bits_addr = readRespArb_io_out_bits_addr; // @[ICache.scala 215:18]
  assign io_read_resp_bits_inst_0 = readRespArb_io_out_bits_inst_0; // @[ICache.scala 215:18]
  assign io_read_resp_bits_inst_1 = readRespArb_io_out_bits_inst_1; // @[ICache.scala 215:18]
  assign io_read_resp_bits_inst_2 = readRespArb_io_out_bits_inst_2; // @[ICache.scala 215:18]
  assign io_read_resp_bits_inst_3 = readRespArb_io_out_bits_inst_3; // @[ICache.scala 215:18]
  assign io_read_resp_bits_size = readRespArb_io_out_bits_size; // @[ICache.scala 215:18]
  assign io_tlbus_req_valid = refillPipe_io_tlbus_req_valid; // @[ICache.scala 66:25]
  assign io_tlbus_req_bits_address = refillPipe_io_tlbus_req_bits_address; // @[ICache.scala 66:25]
  assign io_tlbus_resp_ready = 1'h1; // @[ICache.scala 254:25]
  assign db_clock = clock;
  assign db_reset = reset;
  assign db_io_read_req_valid = s0_latch | s0_full; // @[ICache.scala 88:38]
  assign db_io_read_req_bits_set = _GEN_0[11:5]; // @[Parameters.scala 50:11]
  assign db_io_write_req_valid = refillPipe_io_dataWrite_req_valid; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_set = refillPipe_io_dataWrite_req_bits_set; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_data_0 = refillPipe_io_dataWrite_req_bits_data_0; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_data_1 = refillPipe_io_dataWrite_req_bits_data_1; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_data_2 = refillPipe_io_dataWrite_req_bits_data_2; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_data_3 = refillPipe_io_dataWrite_req_bits_data_3; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_data_4 = refillPipe_io_dataWrite_req_bits_data_4; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_data_5 = refillPipe_io_dataWrite_req_bits_data_5; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_data_6 = refillPipe_io_dataWrite_req_bits_data_6; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_data_7 = refillPipe_io_dataWrite_req_bits_data_7; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_blockMask = refillPipe_io_dataWrite_req_bits_blockMask; // @[ICache.scala 64:33]
  assign db_io_write_req_bits_way = refillPipe_io_dataWrite_req_bits_way; // @[ICache.scala 64:33]
  assign dir_clock = clock;
  assign dir_reset = reset;
  assign dir_io_read_req_valid = s0_latch | s0_full; // @[ICache.scala 91:39]
  assign dir_io_read_req_bits_addr = s0_latch ? io_read_req_bits_addr : s0_req_r_addr; // @[ICache.scala 81:21]
  assign dir_io_write_req_valid = refillPipe_io_dirWrite_req_valid; // @[ICache.scala 65:32]
  assign dir_io_write_req_bits_addr = refillPipe_io_dirWrite_req_bits_addr; // @[ICache.scala 65:32]
  assign dir_io_write_req_bits_way = refillPipe_io_dirWrite_req_bits_way; // @[ICache.scala 65:32]
  assign refillPipe_clock = clock;
  assign refillPipe_reset = reset;
  assign refillPipe_io_req_valid = _s1_resp_valid_T & s1_full & _s1_valid_T_5; // @[ICache.scala 136:64]
  assign refillPipe_io_req_bits_addr = s1_info_req_addr; // @[ICache.scala 137:33]
  assign refillPipe_io_req_bits_chosenWay = s1_info_dirInfo_chosenWay; // @[ICache.scala 138:38]
  assign refillPipe_io_resp_ready = io_read_resp_ready; // @[ICache.scala 252:30]
  assign refillPipe_io_tlbus_req_ready = io_tlbus_req_ready; // @[ICache.scala 66:25]
  assign refillPipe_io_tlbus_resp_valid = io_tlbus_resp_valid; // @[ICache.scala 66:25]
  assign refillPipe_io_tlbus_resp_bits_opcode = io_tlbus_resp_bits_opcode; // @[ICache.scala 66:25]
  assign refillPipe_io_tlbus_resp_bits_data = io_tlbus_resp_bits_data; // @[ICache.scala 66:25]
  assign refillBuffer_clock = clock;
  assign refillBuffer_reset = reset;
  assign refillBuffer_io_write_valid = _refillBuffer_io_write_valid_T & io_tlbus_resp_bits_opcode == 3'h1; // @[ICache.scala 179:55]
  assign refillBuffer_io_write_bits_cacheLineAddr = s2_addr; // @[ICache.scala 181:46]
  assign refillBuffer_io_write_bits_data = io_tlbus_resp_bits_data; // @[ICache.scala 180:37]
  assign readRespArb_io_in_0_valid = _s2_valid_T_1 & s2_full & (_s2_resp_valid_T_2 | s2_refillValid); // @[ICache.scala 193:49]
  assign readRespArb_io_in_0_bits_data = refillPipe_io_resp_bits_data; // @[ICache.scala 192:27 196:23]
  assign readRespArb_io_in_0_bits_addr = s2_addr; // @[ICache.scala 192:27 194:23]
  assign readRespArb_io_in_0_bits_inst_0 = _s2_respRefillInst_T_2[31:0]; // @[ICache.scala 191:133]
  assign readRespArb_io_in_0_bits_inst_1 = _s2_respRefillInst_T_2[63:32]; // @[ICache.scala 191:133]
  assign readRespArb_io_in_0_bits_inst_2 = _s2_respRefillInst_T_2[95:64]; // @[ICache.scala 191:133]
  assign readRespArb_io_in_0_bits_inst_3 = _s2_respRefillInst_T_2[127:96]; // @[ICache.scala 191:133]
  assign readRespArb_io_in_0_bits_size = s2_respMissSize[2:0]; // @[ICache.scala 192:27 195:23]
  assign readRespArb_io_in_1_valid = (s1_info_dirInfo_hit | ~s1_info_dirInfo_hit & s1_bypass) & s1_full & s2_ready; // @[ICache.scala 147:94]
  assign readRespArb_io_in_1_bits_data = s1_bypass ? s1_bypassData : s1_rdHitData; // @[ICache.scala 150:29]
  assign readRespArb_io_in_1_bits_addr = s1_info_req_addr; // @[ICache.scala 146:27 148:23]
  assign readRespArb_io_in_1_bits_inst_0 = s1_bypass ? s1_respBypassInst_0 : s1_respHitInst_0; // @[ICache.scala 152:20]
  assign readRespArb_io_in_1_bits_inst_1 = s1_bypass ? s1_respBypassInst_1 : s1_respHitInst_1; // @[ICache.scala 152:20]
  assign readRespArb_io_in_1_bits_inst_2 = s1_bypass ? s1_respBypassInst_2 : s1_respHitInst_2; // @[ICache.scala 152:20]
  assign readRespArb_io_in_1_bits_inst_3 = s1_bypass ? s1_respBypassInst_3 : s1_respHitInst_3; // @[ICache.scala 152:20]
  assign readRespArb_io_in_1_bits_size = s1_respHitSize[2:0]; // @[ICache.scala 146:27 149:23]
  assign readRespArb_io_out_ready = io_read_resp_ready; // @[ICache.scala 215:18]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 78:26]
      s0_full <= 1'h0; // @[ICache.scala 78:26]
    end else begin
      s0_full <= _GEN_2;
    end
    if (reset) begin // @[ICache.scala 116:26]
      s1_full <= 1'h0; // @[ICache.scala 116:26]
    end else if (io_flush) begin // @[ICache.scala 206:20]
      s1_full <= 1'h0; // @[ICache.scala 207:17]
    end else begin
      s1_full <= _GEN_80;
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_dirInfo_hit <= s0_info_dirInfo_hit; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      if (s0_latch) begin // @[Reg.scala 20:18]
        s1_info_req_addr <= io_read_req_bits_addr; // @[Reg.scala 20:22]
      end else begin
        s1_info_req_addr <= s0_req_r_addr; // @[Reg.scala 19:16]
      end
    end
    if (reset) begin // @[ICache.scala 167:26]
      s2_full <= 1'h0; // @[ICache.scala 167:26]
    end else if (io_flush) begin // @[ICache.scala 206:20]
      s2_full <= 1'h0; // @[ICache.scala 208:17]
    end else begin
      s2_full <= _GEN_111;
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_dirInfo_hit <= s1_info_dirInfo_hit; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_bypass <= s1_bypass; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[ICache.scala 185:33]
      s2_refillValid <= 1'h0; // @[ICache.scala 185:33]
    end else if (s2_refillValid & s1_fire | s2_fire) begin // @[ICache.scala 186:50]
      s2_refillValid <= 1'h0; // @[ICache.scala 186:67]
    end else begin
      s2_refillValid <= _s2_resp_valid_T_3;
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_req_r_addr <= io_read_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_dirInfo_chosenWay <= s0_info_dirInfo_chosenWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_0 <= s0_info_rdData_0_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_1 <= s0_info_rdData_0_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_2 <= s0_info_rdData_0_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_3 <= s0_info_rdData_0_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_4 <= s0_info_rdData_0_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_5 <= s0_info_rdData_0_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_6 <= s0_info_rdData_0_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_7 <= s0_info_rdData_0_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_0 <= s0_info_rdData_1_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_1 <= s0_info_rdData_1_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_2 <= s0_info_rdData_1_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_3 <= s0_info_rdData_1_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_4 <= s0_info_rdData_1_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_5 <= s0_info_rdData_1_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_6 <= s0_info_rdData_1_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_7 <= s0_info_rdData_1_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_0 <= s0_info_rdData_2_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_1 <= s0_info_rdData_2_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_2 <= s0_info_rdData_2_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_3 <= s0_info_rdData_2_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_4 <= s0_info_rdData_2_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_5 <= s0_info_rdData_2_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_6 <= s0_info_rdData_2_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_7 <= s0_info_rdData_2_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_0 <= s0_info_rdData_3_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_1 <= s0_info_rdData_3_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_2 <= s0_info_rdData_3_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_3 <= s0_info_rdData_3_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_4 <= s0_info_rdData_3_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_5 <= s0_info_rdData_3_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_6 <= s0_info_rdData_3_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_7 <= s0_info_rdData_3_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_0 <= s0_info_rdData_4_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_1 <= s0_info_rdData_4_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_2 <= s0_info_rdData_4_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_3 <= s0_info_rdData_4_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_4 <= s0_info_rdData_4_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_5 <= s0_info_rdData_4_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_6 <= s0_info_rdData_4_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_7 <= s0_info_rdData_4_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_0 <= s0_info_rdData_5_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_1 <= s0_info_rdData_5_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_2 <= s0_info_rdData_5_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_3 <= s0_info_rdData_5_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_4 <= s0_info_rdData_5_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_5 <= s0_info_rdData_5_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_6 <= s0_info_rdData_5_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_7 <= s0_info_rdData_5_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_0 <= s0_info_rdData_6_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_1 <= s0_info_rdData_6_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_2 <= s0_info_rdData_6_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_3 <= s0_info_rdData_6_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_4 <= s0_info_rdData_6_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_5 <= s0_info_rdData_6_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_6 <= s0_info_rdData_6_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_7 <= s0_info_rdData_6_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_0 <= s0_info_rdData_7_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_1 <= s0_info_rdData_7_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_2 <= s0_info_rdData_7_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_3 <= s0_info_rdData_7_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_4 <= s0_info_rdData_7_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_5 <= s0_info_rdData_7_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_6 <= s0_info_rdData_7_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_7 <= s0_info_rdData_7_7; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_addr <= s1_info_req_addr; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s1_full = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s1_info_dirInfo_hit = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s1_info_req_addr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  s2_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s2_dirInfo_hit = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s2_bypass = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s2_refillValid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s0_req_r_addr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  s1_info_dirInfo_chosenWay = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  s1_info_rdData_0_0 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  s1_info_rdData_0_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  s1_info_rdData_0_2 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  s1_info_rdData_0_3 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  s1_info_rdData_0_4 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  s1_info_rdData_0_5 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  s1_info_rdData_0_6 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  s1_info_rdData_0_7 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  s1_info_rdData_1_0 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  s1_info_rdData_1_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  s1_info_rdData_1_2 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  s1_info_rdData_1_3 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  s1_info_rdData_1_4 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  s1_info_rdData_1_5 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  s1_info_rdData_1_6 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  s1_info_rdData_1_7 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  s1_info_rdData_2_0 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  s1_info_rdData_2_1 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  s1_info_rdData_2_2 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  s1_info_rdData_2_3 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  s1_info_rdData_2_4 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  s1_info_rdData_2_5 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  s1_info_rdData_2_6 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  s1_info_rdData_2_7 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  s1_info_rdData_3_0 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  s1_info_rdData_3_1 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  s1_info_rdData_3_2 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  s1_info_rdData_3_3 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  s1_info_rdData_3_4 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  s1_info_rdData_3_5 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  s1_info_rdData_3_6 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  s1_info_rdData_3_7 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  s1_info_rdData_4_0 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  s1_info_rdData_4_1 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  s1_info_rdData_4_2 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  s1_info_rdData_4_3 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  s1_info_rdData_4_4 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  s1_info_rdData_4_5 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  s1_info_rdData_4_6 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  s1_info_rdData_4_7 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  s1_info_rdData_5_0 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  s1_info_rdData_5_1 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  s1_info_rdData_5_2 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  s1_info_rdData_5_3 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  s1_info_rdData_5_4 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  s1_info_rdData_5_5 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  s1_info_rdData_5_6 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  s1_info_rdData_5_7 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  s1_info_rdData_6_0 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  s1_info_rdData_6_1 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  s1_info_rdData_6_2 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  s1_info_rdData_6_3 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  s1_info_rdData_6_4 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  s1_info_rdData_6_5 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  s1_info_rdData_6_6 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  s1_info_rdData_6_7 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  s1_info_rdData_7_0 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  s1_info_rdData_7_1 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  s1_info_rdData_7_2 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  s1_info_rdData_7_3 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  s1_info_rdData_7_4 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  s1_info_rdData_7_5 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  s1_info_rdData_7_6 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  s1_info_rdData_7_7 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  s2_addr = _RAND_74[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFile2(
  input         clock,
  input         reset,
  input  [4:0]  io_r_0_addr,
  output [31:0] io_r_0_data,
  input  [4:0]  io_r_1_addr,
  output [31:0] io_r_1_data,
  input  [4:0]  io_r_2_addr,
  output [31:0] io_r_2_data,
  input  [4:0]  io_r_3_addr,
  output [31:0] io_r_3_data,
  input  [4:0]  io_r_4_addr,
  output [31:0] io_r_4_data,
  input  [4:0]  io_r_5_addr,
  output [31:0] io_r_5_data,
  input  [4:0]  io_r_6_addr,
  output [31:0] io_r_6_data,
  input  [4:0]  io_r_7_addr,
  output [31:0] io_r_7_data,
  input  [4:0]  io_w_0_addr,
  input         io_w_0_en,
  input  [31:0] io_w_0_data,
  output [31:0] regState_0_regState_0,
  output [31:0] regState_0_regState_1,
  output [31:0] regState_0_regState_2,
  output [31:0] regState_0_regState_3,
  output [31:0] regState_0_regState_4,
  output [31:0] regState_0_regState_5,
  output [31:0] regState_0_regState_6,
  output [31:0] regState_0_regState_7,
  output [31:0] regState_0_regState_8,
  output [31:0] regState_0_regState_9,
  output [31:0] regState_0_regState_10,
  output [31:0] regState_0_regState_11,
  output [31:0] regState_0_regState_12,
  output [31:0] regState_0_regState_13,
  output [31:0] regState_0_regState_14,
  output [31:0] regState_0_regState_15,
  output [31:0] regState_0_regState_16,
  output [31:0] regState_0_regState_17,
  output [31:0] regState_0_regState_18,
  output [31:0] regState_0_regState_19,
  output [31:0] regState_0_regState_20,
  output [31:0] regState_0_regState_21,
  output [31:0] regState_0_regState_22,
  output [31:0] regState_0_regState_23,
  output [31:0] regState_0_regState_24,
  output [31:0] regState_0_regState_25,
  output [31:0] regState_0_regState_26,
  output [31:0] regState_0_regState_27,
  output [31:0] regState_0_regState_28,
  output [31:0] regState_0_regState_29,
  output [31:0] regState_0_regState_30,
  output [31:0] regState_0_regState_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[RegFile.scala 125:17]
  reg [31:0] regs_1; // @[RegFile.scala 125:17]
  reg [31:0] regs_2; // @[RegFile.scala 125:17]
  reg [31:0] regs_3; // @[RegFile.scala 125:17]
  reg [31:0] regs_4; // @[RegFile.scala 125:17]
  reg [31:0] regs_5; // @[RegFile.scala 125:17]
  reg [31:0] regs_6; // @[RegFile.scala 125:17]
  reg [31:0] regs_7; // @[RegFile.scala 125:17]
  reg [31:0] regs_8; // @[RegFile.scala 125:17]
  reg [31:0] regs_9; // @[RegFile.scala 125:17]
  reg [31:0] regs_10; // @[RegFile.scala 125:17]
  reg [31:0] regs_11; // @[RegFile.scala 125:17]
  reg [31:0] regs_12; // @[RegFile.scala 125:17]
  reg [31:0] regs_13; // @[RegFile.scala 125:17]
  reg [31:0] regs_14; // @[RegFile.scala 125:17]
  reg [31:0] regs_15; // @[RegFile.scala 125:17]
  reg [31:0] regs_16; // @[RegFile.scala 125:17]
  reg [31:0] regs_17; // @[RegFile.scala 125:17]
  reg [31:0] regs_18; // @[RegFile.scala 125:17]
  reg [31:0] regs_19; // @[RegFile.scala 125:17]
  reg [31:0] regs_20; // @[RegFile.scala 125:17]
  reg [31:0] regs_21; // @[RegFile.scala 125:17]
  reg [31:0] regs_22; // @[RegFile.scala 125:17]
  reg [31:0] regs_23; // @[RegFile.scala 125:17]
  reg [31:0] regs_24; // @[RegFile.scala 125:17]
  reg [31:0] regs_25; // @[RegFile.scala 125:17]
  reg [31:0] regs_26; // @[RegFile.scala 125:17]
  reg [31:0] regs_27; // @[RegFile.scala 125:17]
  reg [31:0] regs_28; // @[RegFile.scala 125:17]
  reg [31:0] regs_29; // @[RegFile.scala 125:17]
  reg [31:0] regs_30; // @[RegFile.scala 125:17]
  reg [31:0] regs_31; // @[RegFile.scala 125:17]
  wire [31:0] _GEN_1 = reset ? 32'h0 : regs_1; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_2 = reset ? 32'h0 : regs_2; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_3 = reset ? 32'h0 : regs_3; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_4 = reset ? 32'h0 : regs_4; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_5 = reset ? 32'h0 : regs_5; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_6 = reset ? 32'h0 : regs_6; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_7 = reset ? 32'h0 : regs_7; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_8 = reset ? 32'h0 : regs_8; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_9 = reset ? 32'h0 : regs_9; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_10 = reset ? 32'h0 : regs_10; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_11 = reset ? 32'h0 : regs_11; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_12 = reset ? 32'h0 : regs_12; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_13 = reset ? 32'h0 : regs_13; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_14 = reset ? 32'h0 : regs_14; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_15 = reset ? 32'h0 : regs_15; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_16 = reset ? 32'h0 : regs_16; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_17 = reset ? 32'h0 : regs_17; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_18 = reset ? 32'h0 : regs_18; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_19 = reset ? 32'h0 : regs_19; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_20 = reset ? 32'h0 : regs_20; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_21 = reset ? 32'h0 : regs_21; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_22 = reset ? 32'h0 : regs_22; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_23 = reset ? 32'h0 : regs_23; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_24 = reset ? 32'h0 : regs_24; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_25 = reset ? 32'h0 : regs_25; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_26 = reset ? 32'h0 : regs_26; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_27 = reset ? 32'h0 : regs_27; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_28 = reset ? 32'h0 : regs_28; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_29 = reset ? 32'h0 : regs_29; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_30 = reset ? 32'h0 : regs_30; // @[RegFile.scala 125:17 126:22 128:9]
  wire [31:0] _GEN_31 = reset ? 32'h0 : regs_31; // @[RegFile.scala 125:17 126:22 128:9]
  wire  _writeVec_T_2 = io_w_0_addr != 5'h0; // @[RegFile.scala 152:75]
  wire  _writeVec_T_3 = io_w_0_addr == io_r_0_addr & io_w_0_en & io_w_0_addr != 5'h0; // @[RegFile.scala 152:65]
  wire [3:0] writeVec = {2'h0,1'h0,_writeVec_T_3}; // @[Cat.scala 33:92]
  wire  hasWrite = |writeVec; // @[RegFile.scala 153:29]
  wire [1:0] io_r_0_data_hi = writeVec[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_r_0_data_lo = writeVec[1:0]; // @[OneHot.scala 31:18]
  wire  _io_r_0_data_T = |io_r_0_data_hi; // @[OneHot.scala 32:14]
  wire [1:0] _io_r_0_data_T_1 = io_r_0_data_hi | io_r_0_data_lo; // @[OneHot.scala 32:28]
  wire [1:0] _io_r_0_data_T_3 = {_io_r_0_data_T,_io_r_0_data_T_1[1]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_33 = 2'h1 == _io_r_0_data_T_3 ? 32'h0 : io_w_0_data; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_34 = 2'h2 == _io_r_0_data_T_3 ? 32'h0 : _GEN_33; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_35 = 2'h3 == _io_r_0_data_T_3 ? 32'h0 : _GEN_34; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_36 = regs_0; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_37 = 5'h1 == io_r_0_addr ? regs_1 : regs_0; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_38 = 5'h2 == io_r_0_addr ? regs_2 : _GEN_37; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_39 = 5'h3 == io_r_0_addr ? regs_3 : _GEN_38; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_40 = 5'h4 == io_r_0_addr ? regs_4 : _GEN_39; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_41 = 5'h5 == io_r_0_addr ? regs_5 : _GEN_40; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_42 = 5'h6 == io_r_0_addr ? regs_6 : _GEN_41; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_43 = 5'h7 == io_r_0_addr ? regs_7 : _GEN_42; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_44 = 5'h8 == io_r_0_addr ? regs_8 : _GEN_43; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_45 = 5'h9 == io_r_0_addr ? regs_9 : _GEN_44; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_46 = 5'ha == io_r_0_addr ? regs_10 : _GEN_45; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_47 = 5'hb == io_r_0_addr ? regs_11 : _GEN_46; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_48 = 5'hc == io_r_0_addr ? regs_12 : _GEN_47; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_49 = 5'hd == io_r_0_addr ? regs_13 : _GEN_48; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_50 = 5'he == io_r_0_addr ? regs_14 : _GEN_49; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_51 = 5'hf == io_r_0_addr ? regs_15 : _GEN_50; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_52 = 5'h10 == io_r_0_addr ? regs_16 : _GEN_51; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_53 = 5'h11 == io_r_0_addr ? regs_17 : _GEN_52; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_54 = 5'h12 == io_r_0_addr ? regs_18 : _GEN_53; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_55 = 5'h13 == io_r_0_addr ? regs_19 : _GEN_54; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_56 = 5'h14 == io_r_0_addr ? regs_20 : _GEN_55; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_57 = 5'h15 == io_r_0_addr ? regs_21 : _GEN_56; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_58 = 5'h16 == io_r_0_addr ? regs_22 : _GEN_57; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_59 = 5'h17 == io_r_0_addr ? regs_23 : _GEN_58; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_60 = 5'h18 == io_r_0_addr ? regs_24 : _GEN_59; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_61 = 5'h19 == io_r_0_addr ? regs_25 : _GEN_60; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_62 = 5'h1a == io_r_0_addr ? regs_26 : _GEN_61; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_63 = 5'h1b == io_r_0_addr ? regs_27 : _GEN_62; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_64 = 5'h1c == io_r_0_addr ? regs_28 : _GEN_63; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_65 = 5'h1d == io_r_0_addr ? regs_29 : _GEN_64; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_66 = 5'h1e == io_r_0_addr ? regs_30 : _GEN_65; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_67 = 5'h1f == io_r_0_addr ? regs_31 : _GEN_66; // @[RegFile.scala 158:{16,16}]
  wire  _writeVec_T_19 = io_w_0_addr == io_r_1_addr & io_w_0_en & io_w_0_addr != 5'h0; // @[RegFile.scala 152:65]
  wire [3:0] writeVec_1 = {2'h0,1'h0,_writeVec_T_19}; // @[Cat.scala 33:92]
  wire  hasWrite_1 = |writeVec_1; // @[RegFile.scala 153:29]
  wire [1:0] io_r_1_data_hi = writeVec_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_r_1_data_lo = writeVec_1[1:0]; // @[OneHot.scala 31:18]
  wire  _io_r_1_data_T = |io_r_1_data_hi; // @[OneHot.scala 32:14]
  wire [1:0] _io_r_1_data_T_1 = io_r_1_data_hi | io_r_1_data_lo; // @[OneHot.scala 32:28]
  wire [1:0] _io_r_1_data_T_3 = {_io_r_1_data_T,_io_r_1_data_T_1[1]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_71 = 2'h1 == _io_r_1_data_T_3 ? 32'h0 : io_w_0_data; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_72 = 2'h2 == _io_r_1_data_T_3 ? 32'h0 : _GEN_71; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_73 = 2'h3 == _io_r_1_data_T_3 ? 32'h0 : _GEN_72; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_75 = 5'h1 == io_r_1_addr ? regs_1 : regs_0; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_76 = 5'h2 == io_r_1_addr ? regs_2 : _GEN_75; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_77 = 5'h3 == io_r_1_addr ? regs_3 : _GEN_76; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_78 = 5'h4 == io_r_1_addr ? regs_4 : _GEN_77; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_79 = 5'h5 == io_r_1_addr ? regs_5 : _GEN_78; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_80 = 5'h6 == io_r_1_addr ? regs_6 : _GEN_79; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_81 = 5'h7 == io_r_1_addr ? regs_7 : _GEN_80; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_82 = 5'h8 == io_r_1_addr ? regs_8 : _GEN_81; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_83 = 5'h9 == io_r_1_addr ? regs_9 : _GEN_82; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_84 = 5'ha == io_r_1_addr ? regs_10 : _GEN_83; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_85 = 5'hb == io_r_1_addr ? regs_11 : _GEN_84; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_86 = 5'hc == io_r_1_addr ? regs_12 : _GEN_85; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_87 = 5'hd == io_r_1_addr ? regs_13 : _GEN_86; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_88 = 5'he == io_r_1_addr ? regs_14 : _GEN_87; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_89 = 5'hf == io_r_1_addr ? regs_15 : _GEN_88; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_90 = 5'h10 == io_r_1_addr ? regs_16 : _GEN_89; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_91 = 5'h11 == io_r_1_addr ? regs_17 : _GEN_90; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_92 = 5'h12 == io_r_1_addr ? regs_18 : _GEN_91; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_93 = 5'h13 == io_r_1_addr ? regs_19 : _GEN_92; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_94 = 5'h14 == io_r_1_addr ? regs_20 : _GEN_93; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_95 = 5'h15 == io_r_1_addr ? regs_21 : _GEN_94; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_96 = 5'h16 == io_r_1_addr ? regs_22 : _GEN_95; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_97 = 5'h17 == io_r_1_addr ? regs_23 : _GEN_96; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_98 = 5'h18 == io_r_1_addr ? regs_24 : _GEN_97; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_99 = 5'h19 == io_r_1_addr ? regs_25 : _GEN_98; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_100 = 5'h1a == io_r_1_addr ? regs_26 : _GEN_99; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_101 = 5'h1b == io_r_1_addr ? regs_27 : _GEN_100; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_102 = 5'h1c == io_r_1_addr ? regs_28 : _GEN_101; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_103 = 5'h1d == io_r_1_addr ? regs_29 : _GEN_102; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_104 = 5'h1e == io_r_1_addr ? regs_30 : _GEN_103; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_105 = 5'h1f == io_r_1_addr ? regs_31 : _GEN_104; // @[RegFile.scala 158:{16,16}]
  wire  _writeVec_T_35 = io_w_0_addr == io_r_2_addr & io_w_0_en & io_w_0_addr != 5'h0; // @[RegFile.scala 152:65]
  wire [3:0] writeVec_2 = {2'h0,1'h0,_writeVec_T_35}; // @[Cat.scala 33:92]
  wire  hasWrite_2 = |writeVec_2; // @[RegFile.scala 153:29]
  wire [1:0] io_r_2_data_hi = writeVec_2[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_r_2_data_lo = writeVec_2[1:0]; // @[OneHot.scala 31:18]
  wire  _io_r_2_data_T = |io_r_2_data_hi; // @[OneHot.scala 32:14]
  wire [1:0] _io_r_2_data_T_1 = io_r_2_data_hi | io_r_2_data_lo; // @[OneHot.scala 32:28]
  wire [1:0] _io_r_2_data_T_3 = {_io_r_2_data_T,_io_r_2_data_T_1[1]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_109 = 2'h1 == _io_r_2_data_T_3 ? 32'h0 : io_w_0_data; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_110 = 2'h2 == _io_r_2_data_T_3 ? 32'h0 : _GEN_109; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_111 = 2'h3 == _io_r_2_data_T_3 ? 32'h0 : _GEN_110; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_113 = 5'h1 == io_r_2_addr ? regs_1 : regs_0; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_114 = 5'h2 == io_r_2_addr ? regs_2 : _GEN_113; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_115 = 5'h3 == io_r_2_addr ? regs_3 : _GEN_114; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_116 = 5'h4 == io_r_2_addr ? regs_4 : _GEN_115; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_117 = 5'h5 == io_r_2_addr ? regs_5 : _GEN_116; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_118 = 5'h6 == io_r_2_addr ? regs_6 : _GEN_117; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_119 = 5'h7 == io_r_2_addr ? regs_7 : _GEN_118; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_120 = 5'h8 == io_r_2_addr ? regs_8 : _GEN_119; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_121 = 5'h9 == io_r_2_addr ? regs_9 : _GEN_120; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_122 = 5'ha == io_r_2_addr ? regs_10 : _GEN_121; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_123 = 5'hb == io_r_2_addr ? regs_11 : _GEN_122; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_124 = 5'hc == io_r_2_addr ? regs_12 : _GEN_123; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_125 = 5'hd == io_r_2_addr ? regs_13 : _GEN_124; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_126 = 5'he == io_r_2_addr ? regs_14 : _GEN_125; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_127 = 5'hf == io_r_2_addr ? regs_15 : _GEN_126; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_128 = 5'h10 == io_r_2_addr ? regs_16 : _GEN_127; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_129 = 5'h11 == io_r_2_addr ? regs_17 : _GEN_128; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_130 = 5'h12 == io_r_2_addr ? regs_18 : _GEN_129; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_131 = 5'h13 == io_r_2_addr ? regs_19 : _GEN_130; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_132 = 5'h14 == io_r_2_addr ? regs_20 : _GEN_131; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_133 = 5'h15 == io_r_2_addr ? regs_21 : _GEN_132; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_134 = 5'h16 == io_r_2_addr ? regs_22 : _GEN_133; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_135 = 5'h17 == io_r_2_addr ? regs_23 : _GEN_134; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_136 = 5'h18 == io_r_2_addr ? regs_24 : _GEN_135; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_137 = 5'h19 == io_r_2_addr ? regs_25 : _GEN_136; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_138 = 5'h1a == io_r_2_addr ? regs_26 : _GEN_137; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_139 = 5'h1b == io_r_2_addr ? regs_27 : _GEN_138; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_140 = 5'h1c == io_r_2_addr ? regs_28 : _GEN_139; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_141 = 5'h1d == io_r_2_addr ? regs_29 : _GEN_140; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_142 = 5'h1e == io_r_2_addr ? regs_30 : _GEN_141; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_143 = 5'h1f == io_r_2_addr ? regs_31 : _GEN_142; // @[RegFile.scala 158:{16,16}]
  wire  _writeVec_T_51 = io_w_0_addr == io_r_3_addr & io_w_0_en & io_w_0_addr != 5'h0; // @[RegFile.scala 152:65]
  wire [3:0] writeVec_3 = {2'h0,1'h0,_writeVec_T_51}; // @[Cat.scala 33:92]
  wire  hasWrite_3 = |writeVec_3; // @[RegFile.scala 153:29]
  wire [1:0] io_r_3_data_hi = writeVec_3[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_r_3_data_lo = writeVec_3[1:0]; // @[OneHot.scala 31:18]
  wire  _io_r_3_data_T = |io_r_3_data_hi; // @[OneHot.scala 32:14]
  wire [1:0] _io_r_3_data_T_1 = io_r_3_data_hi | io_r_3_data_lo; // @[OneHot.scala 32:28]
  wire [1:0] _io_r_3_data_T_3 = {_io_r_3_data_T,_io_r_3_data_T_1[1]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_147 = 2'h1 == _io_r_3_data_T_3 ? 32'h0 : io_w_0_data; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_148 = 2'h2 == _io_r_3_data_T_3 ? 32'h0 : _GEN_147; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_149 = 2'h3 == _io_r_3_data_T_3 ? 32'h0 : _GEN_148; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_151 = 5'h1 == io_r_3_addr ? regs_1 : regs_0; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_152 = 5'h2 == io_r_3_addr ? regs_2 : _GEN_151; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_153 = 5'h3 == io_r_3_addr ? regs_3 : _GEN_152; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_154 = 5'h4 == io_r_3_addr ? regs_4 : _GEN_153; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_155 = 5'h5 == io_r_3_addr ? regs_5 : _GEN_154; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_156 = 5'h6 == io_r_3_addr ? regs_6 : _GEN_155; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_157 = 5'h7 == io_r_3_addr ? regs_7 : _GEN_156; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_158 = 5'h8 == io_r_3_addr ? regs_8 : _GEN_157; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_159 = 5'h9 == io_r_3_addr ? regs_9 : _GEN_158; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_160 = 5'ha == io_r_3_addr ? regs_10 : _GEN_159; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_161 = 5'hb == io_r_3_addr ? regs_11 : _GEN_160; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_162 = 5'hc == io_r_3_addr ? regs_12 : _GEN_161; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_163 = 5'hd == io_r_3_addr ? regs_13 : _GEN_162; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_164 = 5'he == io_r_3_addr ? regs_14 : _GEN_163; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_165 = 5'hf == io_r_3_addr ? regs_15 : _GEN_164; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_166 = 5'h10 == io_r_3_addr ? regs_16 : _GEN_165; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_167 = 5'h11 == io_r_3_addr ? regs_17 : _GEN_166; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_168 = 5'h12 == io_r_3_addr ? regs_18 : _GEN_167; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_169 = 5'h13 == io_r_3_addr ? regs_19 : _GEN_168; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_170 = 5'h14 == io_r_3_addr ? regs_20 : _GEN_169; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_171 = 5'h15 == io_r_3_addr ? regs_21 : _GEN_170; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_172 = 5'h16 == io_r_3_addr ? regs_22 : _GEN_171; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_173 = 5'h17 == io_r_3_addr ? regs_23 : _GEN_172; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_174 = 5'h18 == io_r_3_addr ? regs_24 : _GEN_173; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_175 = 5'h19 == io_r_3_addr ? regs_25 : _GEN_174; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_176 = 5'h1a == io_r_3_addr ? regs_26 : _GEN_175; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_177 = 5'h1b == io_r_3_addr ? regs_27 : _GEN_176; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_178 = 5'h1c == io_r_3_addr ? regs_28 : _GEN_177; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_179 = 5'h1d == io_r_3_addr ? regs_29 : _GEN_178; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_180 = 5'h1e == io_r_3_addr ? regs_30 : _GEN_179; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_181 = 5'h1f == io_r_3_addr ? regs_31 : _GEN_180; // @[RegFile.scala 158:{16,16}]
  wire  _writeVec_T_67 = io_w_0_addr == io_r_4_addr & io_w_0_en & io_w_0_addr != 5'h0; // @[RegFile.scala 152:65]
  wire [3:0] writeVec_4 = {2'h0,1'h0,_writeVec_T_67}; // @[Cat.scala 33:92]
  wire  hasWrite_4 = |writeVec_4; // @[RegFile.scala 153:29]
  wire [1:0] io_r_4_data_hi = writeVec_4[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_r_4_data_lo = writeVec_4[1:0]; // @[OneHot.scala 31:18]
  wire  _io_r_4_data_T = |io_r_4_data_hi; // @[OneHot.scala 32:14]
  wire [1:0] _io_r_4_data_T_1 = io_r_4_data_hi | io_r_4_data_lo; // @[OneHot.scala 32:28]
  wire [1:0] _io_r_4_data_T_3 = {_io_r_4_data_T,_io_r_4_data_T_1[1]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_185 = 2'h1 == _io_r_4_data_T_3 ? 32'h0 : io_w_0_data; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_186 = 2'h2 == _io_r_4_data_T_3 ? 32'h0 : _GEN_185; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_187 = 2'h3 == _io_r_4_data_T_3 ? 32'h0 : _GEN_186; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_189 = 5'h1 == io_r_4_addr ? regs_1 : regs_0; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_190 = 5'h2 == io_r_4_addr ? regs_2 : _GEN_189; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_191 = 5'h3 == io_r_4_addr ? regs_3 : _GEN_190; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_192 = 5'h4 == io_r_4_addr ? regs_4 : _GEN_191; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_193 = 5'h5 == io_r_4_addr ? regs_5 : _GEN_192; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_194 = 5'h6 == io_r_4_addr ? regs_6 : _GEN_193; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_195 = 5'h7 == io_r_4_addr ? regs_7 : _GEN_194; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_196 = 5'h8 == io_r_4_addr ? regs_8 : _GEN_195; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_197 = 5'h9 == io_r_4_addr ? regs_9 : _GEN_196; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_198 = 5'ha == io_r_4_addr ? regs_10 : _GEN_197; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_199 = 5'hb == io_r_4_addr ? regs_11 : _GEN_198; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_200 = 5'hc == io_r_4_addr ? regs_12 : _GEN_199; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_201 = 5'hd == io_r_4_addr ? regs_13 : _GEN_200; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_202 = 5'he == io_r_4_addr ? regs_14 : _GEN_201; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_203 = 5'hf == io_r_4_addr ? regs_15 : _GEN_202; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_204 = 5'h10 == io_r_4_addr ? regs_16 : _GEN_203; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_205 = 5'h11 == io_r_4_addr ? regs_17 : _GEN_204; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_206 = 5'h12 == io_r_4_addr ? regs_18 : _GEN_205; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_207 = 5'h13 == io_r_4_addr ? regs_19 : _GEN_206; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_208 = 5'h14 == io_r_4_addr ? regs_20 : _GEN_207; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_209 = 5'h15 == io_r_4_addr ? regs_21 : _GEN_208; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_210 = 5'h16 == io_r_4_addr ? regs_22 : _GEN_209; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_211 = 5'h17 == io_r_4_addr ? regs_23 : _GEN_210; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_212 = 5'h18 == io_r_4_addr ? regs_24 : _GEN_211; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_213 = 5'h19 == io_r_4_addr ? regs_25 : _GEN_212; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_214 = 5'h1a == io_r_4_addr ? regs_26 : _GEN_213; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_215 = 5'h1b == io_r_4_addr ? regs_27 : _GEN_214; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_216 = 5'h1c == io_r_4_addr ? regs_28 : _GEN_215; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_217 = 5'h1d == io_r_4_addr ? regs_29 : _GEN_216; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_218 = 5'h1e == io_r_4_addr ? regs_30 : _GEN_217; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_219 = 5'h1f == io_r_4_addr ? regs_31 : _GEN_218; // @[RegFile.scala 158:{16,16}]
  wire  _writeVec_T_83 = io_w_0_addr == io_r_5_addr & io_w_0_en & io_w_0_addr != 5'h0; // @[RegFile.scala 152:65]
  wire [3:0] writeVec_5 = {2'h0,1'h0,_writeVec_T_83}; // @[Cat.scala 33:92]
  wire  hasWrite_5 = |writeVec_5; // @[RegFile.scala 153:29]
  wire [1:0] io_r_5_data_hi = writeVec_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_r_5_data_lo = writeVec_5[1:0]; // @[OneHot.scala 31:18]
  wire  _io_r_5_data_T = |io_r_5_data_hi; // @[OneHot.scala 32:14]
  wire [1:0] _io_r_5_data_T_1 = io_r_5_data_hi | io_r_5_data_lo; // @[OneHot.scala 32:28]
  wire [1:0] _io_r_5_data_T_3 = {_io_r_5_data_T,_io_r_5_data_T_1[1]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_223 = 2'h1 == _io_r_5_data_T_3 ? 32'h0 : io_w_0_data; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_224 = 2'h2 == _io_r_5_data_T_3 ? 32'h0 : _GEN_223; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_225 = 2'h3 == _io_r_5_data_T_3 ? 32'h0 : _GEN_224; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_227 = 5'h1 == io_r_5_addr ? regs_1 : regs_0; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_228 = 5'h2 == io_r_5_addr ? regs_2 : _GEN_227; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_229 = 5'h3 == io_r_5_addr ? regs_3 : _GEN_228; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_230 = 5'h4 == io_r_5_addr ? regs_4 : _GEN_229; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_231 = 5'h5 == io_r_5_addr ? regs_5 : _GEN_230; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_232 = 5'h6 == io_r_5_addr ? regs_6 : _GEN_231; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_233 = 5'h7 == io_r_5_addr ? regs_7 : _GEN_232; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_234 = 5'h8 == io_r_5_addr ? regs_8 : _GEN_233; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_235 = 5'h9 == io_r_5_addr ? regs_9 : _GEN_234; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_236 = 5'ha == io_r_5_addr ? regs_10 : _GEN_235; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_237 = 5'hb == io_r_5_addr ? regs_11 : _GEN_236; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_238 = 5'hc == io_r_5_addr ? regs_12 : _GEN_237; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_239 = 5'hd == io_r_5_addr ? regs_13 : _GEN_238; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_240 = 5'he == io_r_5_addr ? regs_14 : _GEN_239; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_241 = 5'hf == io_r_5_addr ? regs_15 : _GEN_240; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_242 = 5'h10 == io_r_5_addr ? regs_16 : _GEN_241; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_243 = 5'h11 == io_r_5_addr ? regs_17 : _GEN_242; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_244 = 5'h12 == io_r_5_addr ? regs_18 : _GEN_243; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_245 = 5'h13 == io_r_5_addr ? regs_19 : _GEN_244; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_246 = 5'h14 == io_r_5_addr ? regs_20 : _GEN_245; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_247 = 5'h15 == io_r_5_addr ? regs_21 : _GEN_246; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_248 = 5'h16 == io_r_5_addr ? regs_22 : _GEN_247; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_249 = 5'h17 == io_r_5_addr ? regs_23 : _GEN_248; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_250 = 5'h18 == io_r_5_addr ? regs_24 : _GEN_249; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_251 = 5'h19 == io_r_5_addr ? regs_25 : _GEN_250; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_252 = 5'h1a == io_r_5_addr ? regs_26 : _GEN_251; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_253 = 5'h1b == io_r_5_addr ? regs_27 : _GEN_252; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_254 = 5'h1c == io_r_5_addr ? regs_28 : _GEN_253; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_255 = 5'h1d == io_r_5_addr ? regs_29 : _GEN_254; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_256 = 5'h1e == io_r_5_addr ? regs_30 : _GEN_255; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_257 = 5'h1f == io_r_5_addr ? regs_31 : _GEN_256; // @[RegFile.scala 158:{16,16}]
  wire  _writeVec_T_99 = io_w_0_addr == io_r_6_addr & io_w_0_en & io_w_0_addr != 5'h0; // @[RegFile.scala 152:65]
  wire [3:0] writeVec_6 = {2'h0,1'h0,_writeVec_T_99}; // @[Cat.scala 33:92]
  wire  hasWrite_6 = |writeVec_6; // @[RegFile.scala 153:29]
  wire [1:0] io_r_6_data_hi = writeVec_6[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_r_6_data_lo = writeVec_6[1:0]; // @[OneHot.scala 31:18]
  wire  _io_r_6_data_T = |io_r_6_data_hi; // @[OneHot.scala 32:14]
  wire [1:0] _io_r_6_data_T_1 = io_r_6_data_hi | io_r_6_data_lo; // @[OneHot.scala 32:28]
  wire [1:0] _io_r_6_data_T_3 = {_io_r_6_data_T,_io_r_6_data_T_1[1]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_261 = 2'h1 == _io_r_6_data_T_3 ? 32'h0 : io_w_0_data; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_262 = 2'h2 == _io_r_6_data_T_3 ? 32'h0 : _GEN_261; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_263 = 2'h3 == _io_r_6_data_T_3 ? 32'h0 : _GEN_262; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_265 = 5'h1 == io_r_6_addr ? regs_1 : regs_0; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_266 = 5'h2 == io_r_6_addr ? regs_2 : _GEN_265; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_267 = 5'h3 == io_r_6_addr ? regs_3 : _GEN_266; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_268 = 5'h4 == io_r_6_addr ? regs_4 : _GEN_267; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_269 = 5'h5 == io_r_6_addr ? regs_5 : _GEN_268; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_270 = 5'h6 == io_r_6_addr ? regs_6 : _GEN_269; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_271 = 5'h7 == io_r_6_addr ? regs_7 : _GEN_270; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_272 = 5'h8 == io_r_6_addr ? regs_8 : _GEN_271; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_273 = 5'h9 == io_r_6_addr ? regs_9 : _GEN_272; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_274 = 5'ha == io_r_6_addr ? regs_10 : _GEN_273; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_275 = 5'hb == io_r_6_addr ? regs_11 : _GEN_274; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_276 = 5'hc == io_r_6_addr ? regs_12 : _GEN_275; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_277 = 5'hd == io_r_6_addr ? regs_13 : _GEN_276; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_278 = 5'he == io_r_6_addr ? regs_14 : _GEN_277; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_279 = 5'hf == io_r_6_addr ? regs_15 : _GEN_278; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_280 = 5'h10 == io_r_6_addr ? regs_16 : _GEN_279; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_281 = 5'h11 == io_r_6_addr ? regs_17 : _GEN_280; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_282 = 5'h12 == io_r_6_addr ? regs_18 : _GEN_281; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_283 = 5'h13 == io_r_6_addr ? regs_19 : _GEN_282; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_284 = 5'h14 == io_r_6_addr ? regs_20 : _GEN_283; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_285 = 5'h15 == io_r_6_addr ? regs_21 : _GEN_284; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_286 = 5'h16 == io_r_6_addr ? regs_22 : _GEN_285; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_287 = 5'h17 == io_r_6_addr ? regs_23 : _GEN_286; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_288 = 5'h18 == io_r_6_addr ? regs_24 : _GEN_287; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_289 = 5'h19 == io_r_6_addr ? regs_25 : _GEN_288; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_290 = 5'h1a == io_r_6_addr ? regs_26 : _GEN_289; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_291 = 5'h1b == io_r_6_addr ? regs_27 : _GEN_290; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_292 = 5'h1c == io_r_6_addr ? regs_28 : _GEN_291; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_293 = 5'h1d == io_r_6_addr ? regs_29 : _GEN_292; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_294 = 5'h1e == io_r_6_addr ? regs_30 : _GEN_293; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_295 = 5'h1f == io_r_6_addr ? regs_31 : _GEN_294; // @[RegFile.scala 158:{16,16}]
  wire  _writeVec_T_115 = io_w_0_addr == io_r_7_addr & io_w_0_en & io_w_0_addr != 5'h0; // @[RegFile.scala 152:65]
  wire [3:0] writeVec_7 = {2'h0,1'h0,_writeVec_T_115}; // @[Cat.scala 33:92]
  wire  hasWrite_7 = |writeVec_7; // @[RegFile.scala 153:29]
  wire [1:0] io_r_7_data_hi = writeVec_7[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_r_7_data_lo = writeVec_7[1:0]; // @[OneHot.scala 31:18]
  wire  _io_r_7_data_T = |io_r_7_data_hi; // @[OneHot.scala 32:14]
  wire [1:0] _io_r_7_data_T_1 = io_r_7_data_hi | io_r_7_data_lo; // @[OneHot.scala 32:28]
  wire [1:0] _io_r_7_data_T_3 = {_io_r_7_data_T,_io_r_7_data_T_1[1]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_299 = 2'h1 == _io_r_7_data_T_3 ? 32'h0 : io_w_0_data; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_300 = 2'h2 == _io_r_7_data_T_3 ? 32'h0 : _GEN_299; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_301 = 2'h3 == _io_r_7_data_T_3 ? 32'h0 : _GEN_300; // @[RegFile.scala 156:{16,16}]
  wire [31:0] _GEN_303 = 5'h1 == io_r_7_addr ? regs_1 : regs_0; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_304 = 5'h2 == io_r_7_addr ? regs_2 : _GEN_303; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_305 = 5'h3 == io_r_7_addr ? regs_3 : _GEN_304; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_306 = 5'h4 == io_r_7_addr ? regs_4 : _GEN_305; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_307 = 5'h5 == io_r_7_addr ? regs_5 : _GEN_306; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_308 = 5'h6 == io_r_7_addr ? regs_6 : _GEN_307; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_309 = 5'h7 == io_r_7_addr ? regs_7 : _GEN_308; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_310 = 5'h8 == io_r_7_addr ? regs_8 : _GEN_309; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_311 = 5'h9 == io_r_7_addr ? regs_9 : _GEN_310; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_312 = 5'ha == io_r_7_addr ? regs_10 : _GEN_311; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_313 = 5'hb == io_r_7_addr ? regs_11 : _GEN_312; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_314 = 5'hc == io_r_7_addr ? regs_12 : _GEN_313; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_315 = 5'hd == io_r_7_addr ? regs_13 : _GEN_314; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_316 = 5'he == io_r_7_addr ? regs_14 : _GEN_315; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_317 = 5'hf == io_r_7_addr ? regs_15 : _GEN_316; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_318 = 5'h10 == io_r_7_addr ? regs_16 : _GEN_317; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_319 = 5'h11 == io_r_7_addr ? regs_17 : _GEN_318; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_320 = 5'h12 == io_r_7_addr ? regs_18 : _GEN_319; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_321 = 5'h13 == io_r_7_addr ? regs_19 : _GEN_320; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_322 = 5'h14 == io_r_7_addr ? regs_20 : _GEN_321; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_323 = 5'h15 == io_r_7_addr ? regs_21 : _GEN_322; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_324 = 5'h16 == io_r_7_addr ? regs_22 : _GEN_323; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_325 = 5'h17 == io_r_7_addr ? regs_23 : _GEN_324; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_326 = 5'h18 == io_r_7_addr ? regs_24 : _GEN_325; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_327 = 5'h19 == io_r_7_addr ? regs_25 : _GEN_326; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_328 = 5'h1a == io_r_7_addr ? regs_26 : _GEN_327; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_329 = 5'h1b == io_r_7_addr ? regs_27 : _GEN_328; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_330 = 5'h1c == io_r_7_addr ? regs_28 : _GEN_329; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_331 = 5'h1d == io_r_7_addr ? regs_29 : _GEN_330; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_332 = 5'h1e == io_r_7_addr ? regs_30 : _GEN_331; // @[RegFile.scala 158:{16,16}]
  wire [31:0] _GEN_333 = 5'h1f == io_r_7_addr ? regs_31 : _GEN_332; // @[RegFile.scala 158:{16,16}]
  wire [31:0] regState_regState_0 = regs_0; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_1 = regs_1; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_2 = regs_2; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_3 = regs_3; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_4 = regs_4; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_5 = regs_5; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_6 = regs_6; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_7 = regs_7; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_8 = regs_8; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_9 = regs_9; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_10 = regs_10; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_11 = regs_11; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_12 = regs_12; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_13 = regs_13; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_14 = regs_14; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_15 = regs_15; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_16 = regs_16; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_17 = regs_17; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_18 = regs_18; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_19 = regs_19; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_20 = regs_20; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_21 = regs_21; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_22 = regs_22; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_23 = regs_23; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_24 = regs_24; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_25 = regs_25; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_26 = regs_26; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_27 = regs_27; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_28 = regs_28; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_29 = regs_29; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_30 = regs_30; // @[RegFile.scala 182:22 184:7]
  wire [31:0] regState_regState_31 = regs_31; // @[RegFile.scala 182:22 184:7]
  assign io_r_0_data = hasWrite ? _GEN_35 : _GEN_67; // @[RegFile.scala 155:22 156:16 158:16]
  assign io_r_1_data = hasWrite_1 ? _GEN_73 : _GEN_105; // @[RegFile.scala 155:22 156:16 158:16]
  assign io_r_2_data = hasWrite_2 ? _GEN_111 : _GEN_143; // @[RegFile.scala 155:22 156:16 158:16]
  assign io_r_3_data = hasWrite_3 ? _GEN_149 : _GEN_181; // @[RegFile.scala 155:22 156:16 158:16]
  assign io_r_4_data = hasWrite_4 ? _GEN_187 : _GEN_219; // @[RegFile.scala 155:22 156:16 158:16]
  assign io_r_5_data = hasWrite_5 ? _GEN_225 : _GEN_257; // @[RegFile.scala 155:22 156:16 158:16]
  assign io_r_6_data = hasWrite_6 ? _GEN_263 : _GEN_295; // @[RegFile.scala 155:22 156:16 158:16]
  assign io_r_7_data = hasWrite_7 ? _GEN_301 : _GEN_333; // @[RegFile.scala 155:22 156:16 158:16]
  assign regState_0_regState_0 = _GEN_36;
  assign regState_0_regState_1 = regState_regState_1;
  assign regState_0_regState_2 = regState_regState_2;
  assign regState_0_regState_3 = regState_regState_3;
  assign regState_0_regState_4 = regState_regState_4;
  assign regState_0_regState_5 = regState_regState_5;
  assign regState_0_regState_6 = regState_regState_6;
  assign regState_0_regState_7 = regState_regState_7;
  assign regState_0_regState_8 = regState_regState_8;
  assign regState_0_regState_9 = regState_regState_9;
  assign regState_0_regState_10 = regState_regState_10;
  assign regState_0_regState_11 = regState_regState_11;
  assign regState_0_regState_12 = regState_regState_12;
  assign regState_0_regState_13 = regState_regState_13;
  assign regState_0_regState_14 = regState_regState_14;
  assign regState_0_regState_15 = regState_regState_15;
  assign regState_0_regState_16 = regState_regState_16;
  assign regState_0_regState_17 = regState_regState_17;
  assign regState_0_regState_18 = regState_regState_18;
  assign regState_0_regState_19 = regState_regState_19;
  assign regState_0_regState_20 = regState_regState_20;
  assign regState_0_regState_21 = regState_regState_21;
  assign regState_0_regState_22 = regState_regState_22;
  assign regState_0_regState_23 = regState_regState_23;
  assign regState_0_regState_24 = regState_regState_24;
  assign regState_0_regState_25 = regState_regState_25;
  assign regState_0_regState_26 = regState_regState_26;
  assign regState_0_regState_27 = regState_regState_27;
  assign regState_0_regState_28 = regState_regState_28;
  assign regState_0_regState_29 = regState_regState_29;
  assign regState_0_regState_30 = regState_regState_30;
  assign regState_0_regState_31 = regState_regState_31;
  always @(posedge clock) begin
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h0 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_0 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_0 <= 32'h0; // @[RegFile.scala 133:11]
      end
    end else begin
      regs_0 <= 32'h0; // @[RegFile.scala 133:11]
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h1 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_1 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_1 <= _GEN_1;
      end
    end else begin
      regs_1 <= _GEN_1;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h2 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_2 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_2 <= _GEN_2;
      end
    end else begin
      regs_2 <= _GEN_2;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h3 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_3 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_3 <= _GEN_3;
      end
    end else begin
      regs_3 <= _GEN_3;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h4 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_4 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_4 <= _GEN_4;
      end
    end else begin
      regs_4 <= _GEN_4;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h5 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_5 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_5 <= _GEN_5;
      end
    end else begin
      regs_5 <= _GEN_5;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h6 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_6 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_6 <= _GEN_6;
      end
    end else begin
      regs_6 <= _GEN_6;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h7 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_7 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_7 <= _GEN_7;
      end
    end else begin
      regs_7 <= _GEN_7;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h8 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_8 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_8 <= _GEN_8;
      end
    end else begin
      regs_8 <= _GEN_8;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h9 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_9 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_9 <= _GEN_9;
      end
    end else begin
      regs_9 <= _GEN_9;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'ha == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_10 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_10 <= _GEN_10;
      end
    end else begin
      regs_10 <= _GEN_10;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'hb == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_11 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_11 <= _GEN_11;
      end
    end else begin
      regs_11 <= _GEN_11;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'hc == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_12 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_12 <= _GEN_12;
      end
    end else begin
      regs_12 <= _GEN_12;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'hd == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_13 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_13 <= _GEN_13;
      end
    end else begin
      regs_13 <= _GEN_13;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'he == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_14 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_14 <= _GEN_14;
      end
    end else begin
      regs_14 <= _GEN_14;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'hf == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_15 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_15 <= _GEN_15;
      end
    end else begin
      regs_15 <= _GEN_15;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h10 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_16 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_16 <= _GEN_16;
      end
    end else begin
      regs_16 <= _GEN_16;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h11 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_17 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_17 <= _GEN_17;
      end
    end else begin
      regs_17 <= _GEN_17;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h12 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_18 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_18 <= _GEN_18;
      end
    end else begin
      regs_18 <= _GEN_18;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h13 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_19 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_19 <= _GEN_19;
      end
    end else begin
      regs_19 <= _GEN_19;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h14 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_20 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_20 <= _GEN_20;
      end
    end else begin
      regs_20 <= _GEN_20;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h15 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_21 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_21 <= _GEN_21;
      end
    end else begin
      regs_21 <= _GEN_21;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h16 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_22 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_22 <= _GEN_22;
      end
    end else begin
      regs_22 <= _GEN_22;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h17 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_23 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_23 <= _GEN_23;
      end
    end else begin
      regs_23 <= _GEN_23;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h18 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_24 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_24 <= _GEN_24;
      end
    end else begin
      regs_24 <= _GEN_24;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h19 == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_25 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_25 <= _GEN_25;
      end
    end else begin
      regs_25 <= _GEN_25;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h1a == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_26 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_26 <= _GEN_26;
      end
    end else begin
      regs_26 <= _GEN_26;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h1b == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_27 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_27 <= _GEN_27;
      end
    end else begin
      regs_27 <= _GEN_27;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h1c == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_28 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_28 <= _GEN_28;
      end
    end else begin
      regs_28 <= _GEN_28;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h1d == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_29 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_29 <= _GEN_29;
      end
    end else begin
      regs_29 <= _GEN_29;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h1e == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_30 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_30 <= _GEN_30;
      end
    end else begin
      regs_30 <= _GEN_30;
    end
    if (io_w_0_en & _writeVec_T_2) begin // @[RegFile.scala 173:33]
      if (5'h1f == io_w_0_addr) begin // @[RegFile.scala 174:20]
        regs_31 <= io_w_0_data; // @[RegFile.scala 174:20]
      end else begin
        regs_31 <= _GEN_31;
      end
    end else begin
      regs_31 <= _GEN_31;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(regs_0 == 32'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed: zero reg must be 0 !\n    at RegFile.scala:134 assert(regs(0).asUInt === 0.U, \"zero reg must be 0 !\")\n"
            ); // @[RegFile.scala 134:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(regs_0 == 32'h0) & ~reset) begin
          $fatal; // @[RegFile.scala 134:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ROB(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [4:0]  io_enq_bits_rd,
  input  [3:0]  io_enq_bits_fuValid,
  input  [7:0]  io_enq_bits_fuOp,
  input  [31:0] io_enq_bits_pc,
  input  [31:0] io_enq_bits_inst,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_rdWrEn,
  output [4:0]  io_deq_bits_rd,
  output [31:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_id,
  output [31:0] io_deq_bits_brAddr,
  output        io_deq_bits_brTaken,
  output [31:0] io_deq_bits_excpAddr,
  output        io_deq_bits_excpValid,
  output [31:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_inst,
  input         io_rs_0_valid,
  input  [2:0]  io_rs_0_bits_id,
  input         io_rs_1_valid,
  input  [2:0]  io_rs_1_bits_id,
  input         io_rs_2_valid,
  input  [2:0]  io_rs_2_bits_id,
  input         io_rs_3_valid,
  input  [2:0]  io_rs_3_bits_id,
  output        io_read_0_busy,
  output [1:0]  io_read_0_state,
  output [4:0]  io_read_0_rd,
  output [31:0] io_read_0_data,
  output        io_read_1_busy,
  output [1:0]  io_read_1_state,
  output [4:0]  io_read_1_rd,
  output [31:0] io_read_1_data,
  output        io_read_2_busy,
  output [1:0]  io_read_2_state,
  output [4:0]  io_read_2_rd,
  output [31:0] io_read_2_data,
  output        io_read_3_busy,
  output [1:0]  io_read_3_state,
  output [4:0]  io_read_3_rd,
  output [31:0] io_read_3_data,
  output        io_read_4_busy,
  output [1:0]  io_read_4_state,
  output [4:0]  io_read_4_rd,
  output [31:0] io_read_4_data,
  input         io_fu_0_valid,
  input  [2:0]  io_fu_0_bits_id,
  input  [31:0] io_fu_0_bits_data,
  input         io_fu_1_valid,
  input  [2:0]  io_fu_1_bits_id,
  input  [31:0] io_fu_1_bits_data,
  input  [31:0] io_fu_1_bits_brAddr,
  input         io_fu_1_bits_brTaken,
  input         io_fu_2_valid,
  input  [2:0]  io_fu_2_bits_id,
  input  [31:0] io_fu_2_bits_data,
  input         io_fu_3_valid,
  input  [2:0]  io_fu_3_bits_id,
  input  [31:0] io_fu_3_bits_data,
  input  [31:0] io_fu_3_bits_excpAddr,
  input         io_fu_3_bits_excpValid,
  output [2:0]  io_id,
  output [7:0]  io_regStatus_0_owner,
  output [7:0]  io_regStatus_1_owner,
  output [7:0]  io_regStatus_2_owner,
  output [7:0]  io_regStatus_3_owner,
  output [7:0]  io_regStatus_4_owner,
  output [7:0]  io_regStatus_5_owner,
  output [7:0]  io_regStatus_6_owner,
  output [7:0]  io_regStatus_7_owner,
  output [7:0]  io_regStatus_8_owner,
  output [7:0]  io_regStatus_9_owner,
  output [7:0]  io_regStatus_10_owner,
  output [7:0]  io_regStatus_11_owner,
  output [7:0]  io_regStatus_12_owner,
  output [7:0]  io_regStatus_13_owner,
  output [7:0]  io_regStatus_14_owner,
  output [7:0]  io_regStatus_15_owner,
  output [7:0]  io_regStatus_16_owner,
  output [7:0]  io_regStatus_17_owner,
  output [7:0]  io_regStatus_18_owner,
  output [7:0]  io_regStatus_19_owner,
  output [7:0]  io_regStatus_20_owner,
  output [7:0]  io_regStatus_21_owner,
  output [7:0]  io_regStatus_22_owner,
  output [7:0]  io_regStatus_23_owner,
  output [7:0]  io_regStatus_24_owner,
  output [7:0]  io_regStatus_25_owner,
  output [7:0]  io_regStatus_26_owner,
  output [7:0]  io_regStatus_27_owner,
  output [7:0]  io_regStatus_28_owner,
  output [7:0]  io_regStatus_29_owner,
  output [7:0]  io_regStatus_30_owner,
  output [7:0]  io_regStatus_31_owner,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
`endif // RANDOMIZE_REG_INIT
  reg  entries_0_busy; // @[ROB.scala 118:22]
  reg [1:0] entries_0_state; // @[ROB.scala 118:22]
  reg [4:0] entries_0_rd; // @[ROB.scala 118:22]
  reg [31:0] entries_0_data; // @[ROB.scala 118:22]
  reg [31:0] entries_0_brAddr; // @[ROB.scala 118:22]
  reg  entries_0_brTaken; // @[ROB.scala 118:22]
  reg [31:0] entries_0_excpAddr; // @[ROB.scala 118:22]
  reg  entries_0_excpValid; // @[ROB.scala 118:22]
  reg [31:0] entries_0_pc; // @[ROB.scala 118:22]
  reg [31:0] entries_0_inst; // @[ROB.scala 118:22]
  reg  entries_1_busy; // @[ROB.scala 118:22]
  reg [1:0] entries_1_state; // @[ROB.scala 118:22]
  reg [4:0] entries_1_rd; // @[ROB.scala 118:22]
  reg [31:0] entries_1_data; // @[ROB.scala 118:22]
  reg [31:0] entries_1_brAddr; // @[ROB.scala 118:22]
  reg  entries_1_brTaken; // @[ROB.scala 118:22]
  reg [31:0] entries_1_excpAddr; // @[ROB.scala 118:22]
  reg  entries_1_excpValid; // @[ROB.scala 118:22]
  reg [31:0] entries_1_pc; // @[ROB.scala 118:22]
  reg [31:0] entries_1_inst; // @[ROB.scala 118:22]
  reg  entries_2_busy; // @[ROB.scala 118:22]
  reg [1:0] entries_2_state; // @[ROB.scala 118:22]
  reg [4:0] entries_2_rd; // @[ROB.scala 118:22]
  reg [31:0] entries_2_data; // @[ROB.scala 118:22]
  reg [31:0] entries_2_brAddr; // @[ROB.scala 118:22]
  reg  entries_2_brTaken; // @[ROB.scala 118:22]
  reg [31:0] entries_2_excpAddr; // @[ROB.scala 118:22]
  reg  entries_2_excpValid; // @[ROB.scala 118:22]
  reg [31:0] entries_2_pc; // @[ROB.scala 118:22]
  reg [31:0] entries_2_inst; // @[ROB.scala 118:22]
  reg  entries_3_busy; // @[ROB.scala 118:22]
  reg [1:0] entries_3_state; // @[ROB.scala 118:22]
  reg [4:0] entries_3_rd; // @[ROB.scala 118:22]
  reg [31:0] entries_3_data; // @[ROB.scala 118:22]
  reg [31:0] entries_3_brAddr; // @[ROB.scala 118:22]
  reg  entries_3_brTaken; // @[ROB.scala 118:22]
  reg [31:0] entries_3_excpAddr; // @[ROB.scala 118:22]
  reg  entries_3_excpValid; // @[ROB.scala 118:22]
  reg [31:0] entries_3_pc; // @[ROB.scala 118:22]
  reg [31:0] entries_3_inst; // @[ROB.scala 118:22]
  reg  entries_4_busy; // @[ROB.scala 118:22]
  reg [1:0] entries_4_state; // @[ROB.scala 118:22]
  reg [4:0] entries_4_rd; // @[ROB.scala 118:22]
  reg [31:0] entries_4_data; // @[ROB.scala 118:22]
  reg [31:0] entries_4_brAddr; // @[ROB.scala 118:22]
  reg  entries_4_brTaken; // @[ROB.scala 118:22]
  reg [31:0] entries_4_excpAddr; // @[ROB.scala 118:22]
  reg  entries_4_excpValid; // @[ROB.scala 118:22]
  reg [31:0] entries_4_pc; // @[ROB.scala 118:22]
  reg [31:0] entries_4_inst; // @[ROB.scala 118:22]
  reg [7:0] regResStat_0_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_1_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_2_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_3_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_4_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_5_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_6_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_7_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_8_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_9_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_10_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_11_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_12_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_13_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_14_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_15_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_16_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_17_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_18_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_19_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_20_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_21_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_22_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_23_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_24_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_25_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_26_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_27_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_28_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_29_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_30_owner; // @[ROB.scala 119:25]
  reg [7:0] regResStat_31_owner; // @[ROB.scala 119:25]
  reg [2:0] head; // @[ROB.scala 121:23]
  reg [2:0] tail; // @[ROB.scala 122:23]
  reg [2:0] count; // @[ROB.scala 124:24]
  wire  full = count == 3'h5; // @[ROB.scala 125:22]
  wire [2:0] _io_id_T_1 = tail + 3'h1; // @[ROB.scala 133:19]
  wire  _GEN_1 = 3'h1 == tail ? entries_1_busy : entries_0_busy; // @[ROB.scala 134:{30,30}]
  wire  _GEN_2 = 3'h2 == tail ? entries_2_busy : _GEN_1; // @[ROB.scala 134:{30,30}]
  wire  _GEN_3 = 3'h3 == tail ? entries_3_busy : _GEN_2; // @[ROB.scala 134:{30,30}]
  wire  _GEN_4 = 3'h4 == tail ? entries_4_busy : _GEN_3; // @[ROB.scala 134:{30,30}]
  wire [1:0] _GEN_6 = 3'h1 == head ? entries_1_state : entries_0_state; // @[ROB.scala 135:{41,41}]
  wire [1:0] _GEN_7 = 3'h2 == head ? entries_2_state : _GEN_6; // @[ROB.scala 135:{41,41}]
  wire [1:0] _GEN_8 = 3'h3 == head ? entries_3_state : _GEN_7; // @[ROB.scala 135:{41,41}]
  wire [1:0] _GEN_9 = 3'h4 == head ? entries_4_state : _GEN_8; // @[ROB.scala 135:{41,41}]
  wire  _GEN_11 = 3'h1 == head ? entries_1_busy : entries_0_busy; // @[ROB.scala 135:{52,52}]
  wire  _GEN_12 = 3'h2 == head ? entries_2_busy : _GEN_11; // @[ROB.scala 135:{52,52}]
  wire  _GEN_13 = 3'h3 == head ? entries_3_busy : _GEN_12; // @[ROB.scala 135:{52,52}]
  wire  _GEN_14 = 3'h4 == head ? entries_4_busy : _GEN_13; // @[ROB.scala 135:{52,52}]
  wire [31:0] _GEN_16 = 3'h1 == head ? entries_1_data : entries_0_data; // @[ROB.scala 136:{22,22}]
  wire [31:0] _GEN_17 = 3'h2 == head ? entries_2_data : _GEN_16; // @[ROB.scala 136:{22,22}]
  wire [31:0] _GEN_18 = 3'h3 == head ? entries_3_data : _GEN_17; // @[ROB.scala 136:{22,22}]
  wire [4:0] _GEN_21 = 3'h1 == head ? entries_1_rd : entries_0_rd; // @[ROB.scala 137:{20,20}]
  wire [4:0] _GEN_22 = 3'h2 == head ? entries_2_rd : _GEN_21; // @[ROB.scala 137:{20,20}]
  wire [4:0] _GEN_23 = 3'h3 == head ? entries_3_rd : _GEN_22; // @[ROB.scala 137:{20,20}]
  wire [4:0] _GEN_24 = 3'h4 == head ? entries_4_rd : _GEN_23; // @[ROB.scala 137:{20,20}]
  wire [31:0] _GEN_26 = 3'h1 == head ? entries_1_pc : entries_0_pc; // @[ROB.scala 139:{20,20}]
  wire [31:0] _GEN_27 = 3'h2 == head ? entries_2_pc : _GEN_26; // @[ROB.scala 139:{20,20}]
  wire [31:0] _GEN_28 = 3'h3 == head ? entries_3_pc : _GEN_27; // @[ROB.scala 139:{20,20}]
  wire [31:0] _GEN_31 = 3'h1 == head ? entries_1_inst : entries_0_inst; // @[ROB.scala 140:{22,22}]
  wire [31:0] _GEN_32 = 3'h2 == head ? entries_2_inst : _GEN_31; // @[ROB.scala 140:{22,22}]
  wire [31:0] _GEN_33 = 3'h3 == head ? entries_3_inst : _GEN_32; // @[ROB.scala 140:{22,22}]
  wire [31:0] _GEN_36 = 3'h1 == head ? entries_1_brAddr : entries_0_brAddr; // @[ROB.scala 141:{24,24}]
  wire [31:0] _GEN_37 = 3'h2 == head ? entries_2_brAddr : _GEN_36; // @[ROB.scala 141:{24,24}]
  wire [31:0] _GEN_38 = 3'h3 == head ? entries_3_brAddr : _GEN_37; // @[ROB.scala 141:{24,24}]
  wire  _GEN_41 = 3'h1 == head ? entries_1_brTaken : entries_0_brTaken; // @[ROB.scala 142:{25,25}]
  wire  _GEN_42 = 3'h2 == head ? entries_2_brTaken : _GEN_41; // @[ROB.scala 142:{25,25}]
  wire  _GEN_43 = 3'h3 == head ? entries_3_brTaken : _GEN_42; // @[ROB.scala 142:{25,25}]
  wire [31:0] _GEN_46 = 3'h1 == head ? entries_1_excpAddr : entries_0_excpAddr; // @[ROB.scala 143:{26,26}]
  wire [31:0] _GEN_47 = 3'h2 == head ? entries_2_excpAddr : _GEN_46; // @[ROB.scala 143:{26,26}]
  wire [31:0] _GEN_48 = 3'h3 == head ? entries_3_excpAddr : _GEN_47; // @[ROB.scala 143:{26,26}]
  wire  _GEN_51 = 3'h1 == head ? entries_1_excpValid : entries_0_excpValid; // @[ROB.scala 144:{27,27}]
  wire  _GEN_52 = 3'h2 == head ? entries_2_excpValid : _GEN_51; // @[ROB.scala 144:{27,27}]
  wire  _GEN_53 = 3'h3 == head ? entries_3_excpValid : _GEN_52; // @[ROB.scala 144:{27,27}]
  wire [2:0] _io_deq_bits_id_T_1 = head + 3'h1; // @[ROB.scala 145:28]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_55 = 3'h0 == tail | entries_0_busy; // @[ROB.scala 118:22 149:{28,28}]
  wire  _GEN_56 = 3'h1 == tail | entries_1_busy; // @[ROB.scala 118:22 149:{28,28}]
  wire  _GEN_57 = 3'h2 == tail | entries_2_busy; // @[ROB.scala 118:22 149:{28,28}]
  wire  _GEN_58 = 3'h3 == tail | entries_3_busy; // @[ROB.scala 118:22 149:{28,28}]
  wire  _GEN_59 = 3'h4 == tail | entries_4_busy; // @[ROB.scala 118:22 149:{28,28}]
  wire [1:0] _GEN_60 = 3'h0 == tail ? 2'h0 : entries_0_state; // @[ROB.scala 118:22 150:{29,29}]
  wire [1:0] _GEN_61 = 3'h1 == tail ? 2'h0 : entries_1_state; // @[ROB.scala 118:22 150:{29,29}]
  wire [1:0] _GEN_62 = 3'h2 == tail ? 2'h0 : entries_2_state; // @[ROB.scala 118:22 150:{29,29}]
  wire [1:0] _GEN_63 = 3'h3 == tail ? 2'h0 : entries_3_state; // @[ROB.scala 118:22 150:{29,29}]
  wire [1:0] _GEN_64 = 3'h4 == tail ? 2'h0 : entries_4_state; // @[ROB.scala 118:22 150:{29,29}]
  wire [2:0] _regResStat_owner_T_3 = io_enq_bits_rd == 5'h0 ? 3'h0 : _io_id_T_1; // @[ROB.scala 157:36]
  wire [7:0] _regResStat_io_enq_bits_rd_owner = {{5'd0}, _regResStat_owner_T_3}; // @[ROB.scala 157:{30,30}]
  wire [7:0] _GEN_85 = 5'h0 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_0_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_86 = 5'h1 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_1_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_87 = 5'h2 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_2_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_88 = 5'h3 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_3_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_89 = 5'h4 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_4_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_90 = 5'h5 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_5_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_91 = 5'h6 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_6_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_92 = 5'h7 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_7_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_93 = 5'h8 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_8_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_94 = 5'h9 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_9_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_95 = 5'ha == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_10_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_96 = 5'hb == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_11_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_97 = 5'hc == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_12_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_98 = 5'hd == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_13_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_99 = 5'he == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_14_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_100 = 5'hf == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_15_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_101 = 5'h10 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_16_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_102 = 5'h11 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_17_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_103 = 5'h12 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_18_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_104 = 5'h13 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_19_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_105 = 5'h14 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_20_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_106 = 5'h15 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_21_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_107 = 5'h16 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_22_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_108 = 5'h17 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_23_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_109 = 5'h18 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_24_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_110 = 5'h19 == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_25_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_111 = 5'h1a == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_26_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_112 = 5'h1b == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_27_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_113 = 5'h1c == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_28_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_114 = 5'h1d == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_29_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_115 = 5'h1e == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_30_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire [7:0] _GEN_116 = 5'h1f == io_enq_bits_rd ? _regResStat_io_enq_bits_rd_owner : regResStat_31_owner; // @[ROB.scala 119:25 157:{30,30}]
  wire  _GEN_117 = _T ? _GEN_55 : entries_0_busy; // @[ROB.scala 118:22 148:24]
  wire  _GEN_118 = _T ? _GEN_56 : entries_1_busy; // @[ROB.scala 118:22 148:24]
  wire  _GEN_119 = _T ? _GEN_57 : entries_2_busy; // @[ROB.scala 118:22 148:24]
  wire  _GEN_120 = _T ? _GEN_58 : entries_3_busy; // @[ROB.scala 118:22 148:24]
  wire  _GEN_121 = _T ? _GEN_59 : entries_4_busy; // @[ROB.scala 118:22 148:24]
  wire [1:0] _GEN_122 = _T ? _GEN_60 : entries_0_state; // @[ROB.scala 118:22 148:24]
  wire [1:0] _GEN_123 = _T ? _GEN_61 : entries_1_state; // @[ROB.scala 118:22 148:24]
  wire [1:0] _GEN_124 = _T ? _GEN_62 : entries_2_state; // @[ROB.scala 118:22 148:24]
  wire [1:0] _GEN_125 = _T ? _GEN_63 : entries_3_state; // @[ROB.scala 118:22 148:24]
  wire [1:0] _GEN_126 = _T ? _GEN_64 : entries_4_state; // @[ROB.scala 118:22 148:24]
  wire [7:0] _GEN_142 = _T ? _GEN_85 : regResStat_0_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_143 = _T ? _GEN_86 : regResStat_1_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_144 = _T ? _GEN_87 : regResStat_2_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_145 = _T ? _GEN_88 : regResStat_3_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_146 = _T ? _GEN_89 : regResStat_4_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_147 = _T ? _GEN_90 : regResStat_5_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_148 = _T ? _GEN_91 : regResStat_6_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_149 = _T ? _GEN_92 : regResStat_7_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_150 = _T ? _GEN_93 : regResStat_8_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_151 = _T ? _GEN_94 : regResStat_9_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_152 = _T ? _GEN_95 : regResStat_10_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_153 = _T ? _GEN_96 : regResStat_11_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_154 = _T ? _GEN_97 : regResStat_12_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_155 = _T ? _GEN_98 : regResStat_13_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_156 = _T ? _GEN_99 : regResStat_14_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_157 = _T ? _GEN_100 : regResStat_15_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_158 = _T ? _GEN_101 : regResStat_16_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_159 = _T ? _GEN_102 : regResStat_17_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_160 = _T ? _GEN_103 : regResStat_18_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_161 = _T ? _GEN_104 : regResStat_19_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_162 = _T ? _GEN_105 : regResStat_20_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_163 = _T ? _GEN_106 : regResStat_21_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_164 = _T ? _GEN_107 : regResStat_22_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_165 = _T ? _GEN_108 : regResStat_23_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_166 = _T ? _GEN_109 : regResStat_24_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_167 = _T ? _GEN_110 : regResStat_25_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_168 = _T ? _GEN_111 : regResStat_26_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_169 = _T ? _GEN_112 : regResStat_27_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_170 = _T ? _GEN_113 : regResStat_28_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_171 = _T ? _GEN_114 : regResStat_29_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_172 = _T ? _GEN_115 : regResStat_30_owner; // @[ROB.scala 148:24 119:25]
  wire [7:0] _GEN_173 = _T ? _GEN_116 : regResStat_31_owner; // @[ROB.scala 148:24 119:25]
  wire [1:0] _GEN_180 = 3'h0 == head ? 2'h3 : _GEN_122; // @[ROB.scala 164:{29,29}]
  wire [1:0] _GEN_181 = 3'h1 == head ? 2'h3 : _GEN_123; // @[ROB.scala 164:{29,29}]
  wire [1:0] _GEN_182 = 3'h2 == head ? 2'h3 : _GEN_124; // @[ROB.scala 164:{29,29}]
  wire [1:0] _GEN_183 = 3'h3 == head ? 2'h3 : _GEN_125; // @[ROB.scala 164:{29,29}]
  wire [1:0] _GEN_184 = 3'h4 == head ? 2'h3 : _GEN_126; // @[ROB.scala 164:{29,29}]
  wire  _GEN_185 = 3'h0 == head ? 1'h0 : entries_0_brTaken; // @[ROB.scala 118:22 165:{31,31}]
  wire  _GEN_186 = 3'h1 == head ? 1'h0 : entries_1_brTaken; // @[ROB.scala 118:22 165:{31,31}]
  wire  _GEN_187 = 3'h2 == head ? 1'h0 : entries_2_brTaken; // @[ROB.scala 118:22 165:{31,31}]
  wire  _GEN_188 = 3'h3 == head ? 1'h0 : entries_3_brTaken; // @[ROB.scala 118:22 165:{31,31}]
  wire  _GEN_189 = 3'h4 == head ? 1'h0 : entries_4_brTaken; // @[ROB.scala 118:22 165:{31,31}]
  wire  _GEN_190 = 3'h0 == head ? 1'h0 : entries_0_excpValid; // @[ROB.scala 118:22 166:{33,33}]
  wire  _GEN_191 = 3'h1 == head ? 1'h0 : entries_1_excpValid; // @[ROB.scala 118:22 166:{33,33}]
  wire  _GEN_192 = 3'h2 == head ? 1'h0 : entries_2_excpValid; // @[ROB.scala 118:22 166:{33,33}]
  wire  _GEN_193 = 3'h3 == head ? 1'h0 : entries_3_excpValid; // @[ROB.scala 118:22 166:{33,33}]
  wire  _GEN_194 = 3'h4 == head ? 1'h0 : entries_4_excpValid; // @[ROB.scala 118:22 166:{33,33}]
  wire [7:0] _GEN_196 = 5'h1 == _GEN_24 ? regResStat_1_owner : regResStat_0_owner; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_197 = 5'h2 == _GEN_24 ? regResStat_2_owner : _GEN_196; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_198 = 5'h3 == _GEN_24 ? regResStat_3_owner : _GEN_197; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_199 = 5'h4 == _GEN_24 ? regResStat_4_owner : _GEN_198; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_200 = 5'h5 == _GEN_24 ? regResStat_5_owner : _GEN_199; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_201 = 5'h6 == _GEN_24 ? regResStat_6_owner : _GEN_200; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_202 = 5'h7 == _GEN_24 ? regResStat_7_owner : _GEN_201; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_203 = 5'h8 == _GEN_24 ? regResStat_8_owner : _GEN_202; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_204 = 5'h9 == _GEN_24 ? regResStat_9_owner : _GEN_203; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_205 = 5'ha == _GEN_24 ? regResStat_10_owner : _GEN_204; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_206 = 5'hb == _GEN_24 ? regResStat_11_owner : _GEN_205; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_207 = 5'hc == _GEN_24 ? regResStat_12_owner : _GEN_206; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_208 = 5'hd == _GEN_24 ? regResStat_13_owner : _GEN_207; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_209 = 5'he == _GEN_24 ? regResStat_14_owner : _GEN_208; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_210 = 5'hf == _GEN_24 ? regResStat_15_owner : _GEN_209; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_211 = 5'h10 == _GEN_24 ? regResStat_16_owner : _GEN_210; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_212 = 5'h11 == _GEN_24 ? regResStat_17_owner : _GEN_211; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_213 = 5'h12 == _GEN_24 ? regResStat_18_owner : _GEN_212; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_214 = 5'h13 == _GEN_24 ? regResStat_19_owner : _GEN_213; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_215 = 5'h14 == _GEN_24 ? regResStat_20_owner : _GEN_214; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_216 = 5'h15 == _GEN_24 ? regResStat_21_owner : _GEN_215; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_217 = 5'h16 == _GEN_24 ? regResStat_22_owner : _GEN_216; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_218 = 5'h17 == _GEN_24 ? regResStat_23_owner : _GEN_217; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_219 = 5'h18 == _GEN_24 ? regResStat_24_owner : _GEN_218; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_220 = 5'h19 == _GEN_24 ? regResStat_25_owner : _GEN_219; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_221 = 5'h1a == _GEN_24 ? regResStat_26_owner : _GEN_220; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_222 = 5'h1b == _GEN_24 ? regResStat_27_owner : _GEN_221; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_223 = 5'h1c == _GEN_24 ? regResStat_28_owner : _GEN_222; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_224 = 5'h1d == _GEN_24 ? regResStat_29_owner : _GEN_223; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_225 = 5'h1e == _GEN_24 ? regResStat_30_owner : _GEN_224; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_226 = 5'h1f == _GEN_24 ? regResStat_31_owner : _GEN_225; // @[ROB.scala 169:{43,43}]
  wire [7:0] _GEN_672 = {{5'd0}, _io_deq_bits_id_T_1}; // @[ROB.scala 169:43]
  wire [1:0] _GEN_296 = io_deq_valid ? _GEN_180 : _GEN_122; // @[ROB.scala 162:24]
  wire [1:0] _GEN_297 = io_deq_valid ? _GEN_181 : _GEN_123; // @[ROB.scala 162:24]
  wire [1:0] _GEN_298 = io_deq_valid ? _GEN_182 : _GEN_124; // @[ROB.scala 162:24]
  wire [1:0] _GEN_299 = io_deq_valid ? _GEN_183 : _GEN_125; // @[ROB.scala 162:24]
  wire [1:0] _GEN_300 = io_deq_valid ? _GEN_184 : _GEN_126; // @[ROB.scala 162:24]
  wire  _GEN_301 = io_deq_valid ? _GEN_185 : entries_0_brTaken; // @[ROB.scala 118:22 162:24]
  wire  _GEN_302 = io_deq_valid ? _GEN_186 : entries_1_brTaken; // @[ROB.scala 118:22 162:24]
  wire  _GEN_303 = io_deq_valid ? _GEN_187 : entries_2_brTaken; // @[ROB.scala 118:22 162:24]
  wire  _GEN_304 = io_deq_valid ? _GEN_188 : entries_3_brTaken; // @[ROB.scala 118:22 162:24]
  wire  _GEN_305 = io_deq_valid ? _GEN_189 : entries_4_brTaken; // @[ROB.scala 118:22 162:24]
  wire  _GEN_306 = io_deq_valid ? _GEN_190 : entries_0_excpValid; // @[ROB.scala 118:22 162:24]
  wire  _GEN_307 = io_deq_valid ? _GEN_191 : entries_1_excpValid; // @[ROB.scala 118:22 162:24]
  wire  _GEN_308 = io_deq_valid ? _GEN_192 : entries_2_excpValid; // @[ROB.scala 118:22 162:24]
  wire  _GEN_309 = io_deq_valid ? _GEN_193 : entries_3_excpValid; // @[ROB.scala 118:22 162:24]
  wire  _GEN_310 = io_deq_valid ? _GEN_194 : entries_4_excpValid; // @[ROB.scala 118:22 162:24]
  wire [2:0] _count_T_1 = count + 3'h1; // @[ROB.scala 178:28]
  wire [2:0] _GEN_344 = _T ? _count_T_1 : count; // @[ROB.scala 177:27 178:19 124:24]
  wire [2:0] _count_T_3 = count - 3'h1; // @[ROB.scala 181:28]
  wire [2:0] _T_17 = io_fu_0_bits_id - 3'h1; // @[ROB.scala 187:31]
  wire [31:0] _GEN_347 = 3'h0 == _T_17 ? io_fu_0_bits_data : entries_0_data; // @[ROB.scala 118:22 187:{43,43}]
  wire [31:0] _GEN_348 = 3'h1 == _T_17 ? io_fu_0_bits_data : entries_1_data; // @[ROB.scala 118:22 187:{43,43}]
  wire [31:0] _GEN_349 = 3'h2 == _T_17 ? io_fu_0_bits_data : entries_2_data; // @[ROB.scala 118:22 187:{43,43}]
  wire [31:0] _GEN_350 = 3'h3 == _T_17 ? io_fu_0_bits_data : entries_3_data; // @[ROB.scala 118:22 187:{43,43}]
  wire [31:0] _GEN_351 = 3'h4 == _T_17 ? io_fu_0_bits_data : entries_4_data; // @[ROB.scala 118:22 187:{43,43}]
  wire [1:0] _GEN_352 = 3'h0 == _T_17 ? 2'h2 : _GEN_296; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_353 = 3'h1 == _T_17 ? 2'h2 : _GEN_297; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_354 = 3'h2 == _T_17 ? 2'h2 : _GEN_298; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_355 = 3'h3 == _T_17 ? 2'h2 : _GEN_299; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_356 = 3'h4 == _T_17 ? 2'h2 : _GEN_300; // @[ROB.scala 188:{44,44}]
  wire [31:0] _GEN_357 = 3'h0 == _T_17 ? 32'h0 : entries_0_brAddr; // @[ROB.scala 118:22 189:{45,45}]
  wire [31:0] _GEN_358 = 3'h1 == _T_17 ? 32'h0 : entries_1_brAddr; // @[ROB.scala 118:22 189:{45,45}]
  wire [31:0] _GEN_359 = 3'h2 == _T_17 ? 32'h0 : entries_2_brAddr; // @[ROB.scala 118:22 189:{45,45}]
  wire [31:0] _GEN_360 = 3'h3 == _T_17 ? 32'h0 : entries_3_brAddr; // @[ROB.scala 118:22 189:{45,45}]
  wire [31:0] _GEN_361 = 3'h4 == _T_17 ? 32'h0 : entries_4_brAddr; // @[ROB.scala 118:22 189:{45,45}]
  wire  _GEN_362 = 3'h0 == _T_17 ? 1'h0 : _GEN_301; // @[ROB.scala 190:{46,46}]
  wire  _GEN_363 = 3'h1 == _T_17 ? 1'h0 : _GEN_302; // @[ROB.scala 190:{46,46}]
  wire  _GEN_364 = 3'h2 == _T_17 ? 1'h0 : _GEN_303; // @[ROB.scala 190:{46,46}]
  wire  _GEN_365 = 3'h3 == _T_17 ? 1'h0 : _GEN_304; // @[ROB.scala 190:{46,46}]
  wire  _GEN_366 = 3'h4 == _T_17 ? 1'h0 : _GEN_305; // @[ROB.scala 190:{46,46}]
  wire [31:0] _GEN_367 = 3'h0 == _T_17 ? 32'h0 : entries_0_excpAddr; // @[ROB.scala 118:22 191:{47,47}]
  wire [31:0] _GEN_368 = 3'h1 == _T_17 ? 32'h0 : entries_1_excpAddr; // @[ROB.scala 118:22 191:{47,47}]
  wire [31:0] _GEN_369 = 3'h2 == _T_17 ? 32'h0 : entries_2_excpAddr; // @[ROB.scala 118:22 191:{47,47}]
  wire [31:0] _GEN_370 = 3'h3 == _T_17 ? 32'h0 : entries_3_excpAddr; // @[ROB.scala 118:22 191:{47,47}]
  wire [31:0] _GEN_371 = 3'h4 == _T_17 ? 32'h0 : entries_4_excpAddr; // @[ROB.scala 118:22 191:{47,47}]
  wire  _GEN_372 = 3'h0 == _T_17 ? 1'h0 : _GEN_306; // @[ROB.scala 192:{48,48}]
  wire  _GEN_373 = 3'h1 == _T_17 ? 1'h0 : _GEN_307; // @[ROB.scala 192:{48,48}]
  wire  _GEN_374 = 3'h2 == _T_17 ? 1'h0 : _GEN_308; // @[ROB.scala 192:{48,48}]
  wire  _GEN_375 = 3'h3 == _T_17 ? 1'h0 : _GEN_309; // @[ROB.scala 192:{48,48}]
  wire  _GEN_376 = 3'h4 == _T_17 ? 1'h0 : _GEN_310; // @[ROB.scala 192:{48,48}]
  wire [31:0] _GEN_377 = io_fu_0_valid ? _GEN_347 : entries_0_data; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_378 = io_fu_0_valid ? _GEN_348 : entries_1_data; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_379 = io_fu_0_valid ? _GEN_349 : entries_2_data; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_380 = io_fu_0_valid ? _GEN_350 : entries_3_data; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_381 = io_fu_0_valid ? _GEN_351 : entries_4_data; // @[ROB.scala 118:22 186:23]
  wire [1:0] _GEN_382 = io_fu_0_valid ? _GEN_352 : _GEN_296; // @[ROB.scala 186:23]
  wire [1:0] _GEN_383 = io_fu_0_valid ? _GEN_353 : _GEN_297; // @[ROB.scala 186:23]
  wire [1:0] _GEN_384 = io_fu_0_valid ? _GEN_354 : _GEN_298; // @[ROB.scala 186:23]
  wire [1:0] _GEN_385 = io_fu_0_valid ? _GEN_355 : _GEN_299; // @[ROB.scala 186:23]
  wire [1:0] _GEN_386 = io_fu_0_valid ? _GEN_356 : _GEN_300; // @[ROB.scala 186:23]
  wire [31:0] _GEN_387 = io_fu_0_valid ? _GEN_357 : entries_0_brAddr; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_388 = io_fu_0_valid ? _GEN_358 : entries_1_brAddr; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_389 = io_fu_0_valid ? _GEN_359 : entries_2_brAddr; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_390 = io_fu_0_valid ? _GEN_360 : entries_3_brAddr; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_391 = io_fu_0_valid ? _GEN_361 : entries_4_brAddr; // @[ROB.scala 118:22 186:23]
  wire  _GEN_392 = io_fu_0_valid ? _GEN_362 : _GEN_301; // @[ROB.scala 186:23]
  wire  _GEN_393 = io_fu_0_valid ? _GEN_363 : _GEN_302; // @[ROB.scala 186:23]
  wire  _GEN_394 = io_fu_0_valid ? _GEN_364 : _GEN_303; // @[ROB.scala 186:23]
  wire  _GEN_395 = io_fu_0_valid ? _GEN_365 : _GEN_304; // @[ROB.scala 186:23]
  wire  _GEN_396 = io_fu_0_valid ? _GEN_366 : _GEN_305; // @[ROB.scala 186:23]
  wire [31:0] _GEN_397 = io_fu_0_valid ? _GEN_367 : entries_0_excpAddr; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_398 = io_fu_0_valid ? _GEN_368 : entries_1_excpAddr; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_399 = io_fu_0_valid ? _GEN_369 : entries_2_excpAddr; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_400 = io_fu_0_valid ? _GEN_370 : entries_3_excpAddr; // @[ROB.scala 118:22 186:23]
  wire [31:0] _GEN_401 = io_fu_0_valid ? _GEN_371 : entries_4_excpAddr; // @[ROB.scala 118:22 186:23]
  wire  _GEN_402 = io_fu_0_valid ? _GEN_372 : _GEN_306; // @[ROB.scala 186:23]
  wire  _GEN_403 = io_fu_0_valid ? _GEN_373 : _GEN_307; // @[ROB.scala 186:23]
  wire  _GEN_404 = io_fu_0_valid ? _GEN_374 : _GEN_308; // @[ROB.scala 186:23]
  wire  _GEN_405 = io_fu_0_valid ? _GEN_375 : _GEN_309; // @[ROB.scala 186:23]
  wire  _GEN_406 = io_fu_0_valid ? _GEN_376 : _GEN_310; // @[ROB.scala 186:23]
  wire [2:0] _T_29 = io_fu_1_bits_id - 3'h1; // @[ROB.scala 187:31]
  wire [31:0] _GEN_407 = 3'h0 == _T_29 ? io_fu_1_bits_data : _GEN_377; // @[ROB.scala 187:{43,43}]
  wire [31:0] _GEN_408 = 3'h1 == _T_29 ? io_fu_1_bits_data : _GEN_378; // @[ROB.scala 187:{43,43}]
  wire [31:0] _GEN_409 = 3'h2 == _T_29 ? io_fu_1_bits_data : _GEN_379; // @[ROB.scala 187:{43,43}]
  wire [31:0] _GEN_410 = 3'h3 == _T_29 ? io_fu_1_bits_data : _GEN_380; // @[ROB.scala 187:{43,43}]
  wire [31:0] _GEN_411 = 3'h4 == _T_29 ? io_fu_1_bits_data : _GEN_381; // @[ROB.scala 187:{43,43}]
  wire [1:0] _GEN_412 = 3'h0 == _T_29 ? 2'h2 : _GEN_382; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_413 = 3'h1 == _T_29 ? 2'h2 : _GEN_383; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_414 = 3'h2 == _T_29 ? 2'h2 : _GEN_384; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_415 = 3'h3 == _T_29 ? 2'h2 : _GEN_385; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_416 = 3'h4 == _T_29 ? 2'h2 : _GEN_386; // @[ROB.scala 188:{44,44}]
  wire [31:0] _GEN_417 = 3'h0 == _T_29 ? io_fu_1_bits_brAddr : _GEN_387; // @[ROB.scala 189:{45,45}]
  wire [31:0] _GEN_418 = 3'h1 == _T_29 ? io_fu_1_bits_brAddr : _GEN_388; // @[ROB.scala 189:{45,45}]
  wire [31:0] _GEN_419 = 3'h2 == _T_29 ? io_fu_1_bits_brAddr : _GEN_389; // @[ROB.scala 189:{45,45}]
  wire [31:0] _GEN_420 = 3'h3 == _T_29 ? io_fu_1_bits_brAddr : _GEN_390; // @[ROB.scala 189:{45,45}]
  wire [31:0] _GEN_421 = 3'h4 == _T_29 ? io_fu_1_bits_brAddr : _GEN_391; // @[ROB.scala 189:{45,45}]
  wire  _GEN_422 = 3'h0 == _T_29 ? io_fu_1_bits_brTaken : _GEN_392; // @[ROB.scala 190:{46,46}]
  wire  _GEN_423 = 3'h1 == _T_29 ? io_fu_1_bits_brTaken : _GEN_393; // @[ROB.scala 190:{46,46}]
  wire  _GEN_424 = 3'h2 == _T_29 ? io_fu_1_bits_brTaken : _GEN_394; // @[ROB.scala 190:{46,46}]
  wire  _GEN_425 = 3'h3 == _T_29 ? io_fu_1_bits_brTaken : _GEN_395; // @[ROB.scala 190:{46,46}]
  wire  _GEN_426 = 3'h4 == _T_29 ? io_fu_1_bits_brTaken : _GEN_396; // @[ROB.scala 190:{46,46}]
  wire [31:0] _GEN_427 = 3'h0 == _T_29 ? 32'h0 : _GEN_397; // @[ROB.scala 191:{47,47}]
  wire [31:0] _GEN_428 = 3'h1 == _T_29 ? 32'h0 : _GEN_398; // @[ROB.scala 191:{47,47}]
  wire [31:0] _GEN_429 = 3'h2 == _T_29 ? 32'h0 : _GEN_399; // @[ROB.scala 191:{47,47}]
  wire [31:0] _GEN_430 = 3'h3 == _T_29 ? 32'h0 : _GEN_400; // @[ROB.scala 191:{47,47}]
  wire [31:0] _GEN_431 = 3'h4 == _T_29 ? 32'h0 : _GEN_401; // @[ROB.scala 191:{47,47}]
  wire  _GEN_432 = 3'h0 == _T_29 ? 1'h0 : _GEN_402; // @[ROB.scala 192:{48,48}]
  wire  _GEN_433 = 3'h1 == _T_29 ? 1'h0 : _GEN_403; // @[ROB.scala 192:{48,48}]
  wire  _GEN_434 = 3'h2 == _T_29 ? 1'h0 : _GEN_404; // @[ROB.scala 192:{48,48}]
  wire  _GEN_435 = 3'h3 == _T_29 ? 1'h0 : _GEN_405; // @[ROB.scala 192:{48,48}]
  wire  _GEN_436 = 3'h4 == _T_29 ? 1'h0 : _GEN_406; // @[ROB.scala 192:{48,48}]
  wire [31:0] _GEN_437 = io_fu_1_valid ? _GEN_407 : _GEN_377; // @[ROB.scala 186:23]
  wire [31:0] _GEN_438 = io_fu_1_valid ? _GEN_408 : _GEN_378; // @[ROB.scala 186:23]
  wire [31:0] _GEN_439 = io_fu_1_valid ? _GEN_409 : _GEN_379; // @[ROB.scala 186:23]
  wire [31:0] _GEN_440 = io_fu_1_valid ? _GEN_410 : _GEN_380; // @[ROB.scala 186:23]
  wire [31:0] _GEN_441 = io_fu_1_valid ? _GEN_411 : _GEN_381; // @[ROB.scala 186:23]
  wire [1:0] _GEN_442 = io_fu_1_valid ? _GEN_412 : _GEN_382; // @[ROB.scala 186:23]
  wire [1:0] _GEN_443 = io_fu_1_valid ? _GEN_413 : _GEN_383; // @[ROB.scala 186:23]
  wire [1:0] _GEN_444 = io_fu_1_valid ? _GEN_414 : _GEN_384; // @[ROB.scala 186:23]
  wire [1:0] _GEN_445 = io_fu_1_valid ? _GEN_415 : _GEN_385; // @[ROB.scala 186:23]
  wire [1:0] _GEN_446 = io_fu_1_valid ? _GEN_416 : _GEN_386; // @[ROB.scala 186:23]
  wire [31:0] _GEN_447 = io_fu_1_valid ? _GEN_417 : _GEN_387; // @[ROB.scala 186:23]
  wire [31:0] _GEN_448 = io_fu_1_valid ? _GEN_418 : _GEN_388; // @[ROB.scala 186:23]
  wire [31:0] _GEN_449 = io_fu_1_valid ? _GEN_419 : _GEN_389; // @[ROB.scala 186:23]
  wire [31:0] _GEN_450 = io_fu_1_valid ? _GEN_420 : _GEN_390; // @[ROB.scala 186:23]
  wire [31:0] _GEN_451 = io_fu_1_valid ? _GEN_421 : _GEN_391; // @[ROB.scala 186:23]
  wire  _GEN_452 = io_fu_1_valid ? _GEN_422 : _GEN_392; // @[ROB.scala 186:23]
  wire  _GEN_453 = io_fu_1_valid ? _GEN_423 : _GEN_393; // @[ROB.scala 186:23]
  wire  _GEN_454 = io_fu_1_valid ? _GEN_424 : _GEN_394; // @[ROB.scala 186:23]
  wire  _GEN_455 = io_fu_1_valid ? _GEN_425 : _GEN_395; // @[ROB.scala 186:23]
  wire  _GEN_456 = io_fu_1_valid ? _GEN_426 : _GEN_396; // @[ROB.scala 186:23]
  wire [31:0] _GEN_457 = io_fu_1_valid ? _GEN_427 : _GEN_397; // @[ROB.scala 186:23]
  wire [31:0] _GEN_458 = io_fu_1_valid ? _GEN_428 : _GEN_398; // @[ROB.scala 186:23]
  wire [31:0] _GEN_459 = io_fu_1_valid ? _GEN_429 : _GEN_399; // @[ROB.scala 186:23]
  wire [31:0] _GEN_460 = io_fu_1_valid ? _GEN_430 : _GEN_400; // @[ROB.scala 186:23]
  wire [31:0] _GEN_461 = io_fu_1_valid ? _GEN_431 : _GEN_401; // @[ROB.scala 186:23]
  wire  _GEN_462 = io_fu_1_valid ? _GEN_432 : _GEN_402; // @[ROB.scala 186:23]
  wire  _GEN_463 = io_fu_1_valid ? _GEN_433 : _GEN_403; // @[ROB.scala 186:23]
  wire  _GEN_464 = io_fu_1_valid ? _GEN_434 : _GEN_404; // @[ROB.scala 186:23]
  wire  _GEN_465 = io_fu_1_valid ? _GEN_435 : _GEN_405; // @[ROB.scala 186:23]
  wire  _GEN_466 = io_fu_1_valid ? _GEN_436 : _GEN_406; // @[ROB.scala 186:23]
  wire [2:0] _T_41 = io_fu_2_bits_id - 3'h1; // @[ROB.scala 187:31]
  wire [31:0] _GEN_467 = 3'h0 == _T_41 ? io_fu_2_bits_data : _GEN_437; // @[ROB.scala 187:{43,43}]
  wire [31:0] _GEN_468 = 3'h1 == _T_41 ? io_fu_2_bits_data : _GEN_438; // @[ROB.scala 187:{43,43}]
  wire [31:0] _GEN_469 = 3'h2 == _T_41 ? io_fu_2_bits_data : _GEN_439; // @[ROB.scala 187:{43,43}]
  wire [31:0] _GEN_470 = 3'h3 == _T_41 ? io_fu_2_bits_data : _GEN_440; // @[ROB.scala 187:{43,43}]
  wire [31:0] _GEN_471 = 3'h4 == _T_41 ? io_fu_2_bits_data : _GEN_441; // @[ROB.scala 187:{43,43}]
  wire [1:0] _GEN_472 = 3'h0 == _T_41 ? 2'h2 : _GEN_442; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_473 = 3'h1 == _T_41 ? 2'h2 : _GEN_443; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_474 = 3'h2 == _T_41 ? 2'h2 : _GEN_444; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_475 = 3'h3 == _T_41 ? 2'h2 : _GEN_445; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_476 = 3'h4 == _T_41 ? 2'h2 : _GEN_446; // @[ROB.scala 188:{44,44}]
  wire [31:0] _GEN_477 = 3'h0 == _T_41 ? 32'h0 : _GEN_447; // @[ROB.scala 189:{45,45}]
  wire [31:0] _GEN_478 = 3'h1 == _T_41 ? 32'h0 : _GEN_448; // @[ROB.scala 189:{45,45}]
  wire [31:0] _GEN_479 = 3'h2 == _T_41 ? 32'h0 : _GEN_449; // @[ROB.scala 189:{45,45}]
  wire [31:0] _GEN_480 = 3'h3 == _T_41 ? 32'h0 : _GEN_450; // @[ROB.scala 189:{45,45}]
  wire [31:0] _GEN_481 = 3'h4 == _T_41 ? 32'h0 : _GEN_451; // @[ROB.scala 189:{45,45}]
  wire  _GEN_482 = 3'h0 == _T_41 ? 1'h0 : _GEN_452; // @[ROB.scala 190:{46,46}]
  wire  _GEN_483 = 3'h1 == _T_41 ? 1'h0 : _GEN_453; // @[ROB.scala 190:{46,46}]
  wire  _GEN_484 = 3'h2 == _T_41 ? 1'h0 : _GEN_454; // @[ROB.scala 190:{46,46}]
  wire  _GEN_485 = 3'h3 == _T_41 ? 1'h0 : _GEN_455; // @[ROB.scala 190:{46,46}]
  wire  _GEN_486 = 3'h4 == _T_41 ? 1'h0 : _GEN_456; // @[ROB.scala 190:{46,46}]
  wire [31:0] _GEN_487 = 3'h0 == _T_41 ? 32'h0 : _GEN_457; // @[ROB.scala 191:{47,47}]
  wire [31:0] _GEN_488 = 3'h1 == _T_41 ? 32'h0 : _GEN_458; // @[ROB.scala 191:{47,47}]
  wire [31:0] _GEN_489 = 3'h2 == _T_41 ? 32'h0 : _GEN_459; // @[ROB.scala 191:{47,47}]
  wire [31:0] _GEN_490 = 3'h3 == _T_41 ? 32'h0 : _GEN_460; // @[ROB.scala 191:{47,47}]
  wire [31:0] _GEN_491 = 3'h4 == _T_41 ? 32'h0 : _GEN_461; // @[ROB.scala 191:{47,47}]
  wire  _GEN_492 = 3'h0 == _T_41 ? 1'h0 : _GEN_462; // @[ROB.scala 192:{48,48}]
  wire  _GEN_493 = 3'h1 == _T_41 ? 1'h0 : _GEN_463; // @[ROB.scala 192:{48,48}]
  wire  _GEN_494 = 3'h2 == _T_41 ? 1'h0 : _GEN_464; // @[ROB.scala 192:{48,48}]
  wire  _GEN_495 = 3'h3 == _T_41 ? 1'h0 : _GEN_465; // @[ROB.scala 192:{48,48}]
  wire  _GEN_496 = 3'h4 == _T_41 ? 1'h0 : _GEN_466; // @[ROB.scala 192:{48,48}]
  wire [31:0] _GEN_497 = io_fu_2_valid ? _GEN_467 : _GEN_437; // @[ROB.scala 186:23]
  wire [31:0] _GEN_498 = io_fu_2_valid ? _GEN_468 : _GEN_438; // @[ROB.scala 186:23]
  wire [31:0] _GEN_499 = io_fu_2_valid ? _GEN_469 : _GEN_439; // @[ROB.scala 186:23]
  wire [31:0] _GEN_500 = io_fu_2_valid ? _GEN_470 : _GEN_440; // @[ROB.scala 186:23]
  wire [31:0] _GEN_501 = io_fu_2_valid ? _GEN_471 : _GEN_441; // @[ROB.scala 186:23]
  wire [1:0] _GEN_502 = io_fu_2_valid ? _GEN_472 : _GEN_442; // @[ROB.scala 186:23]
  wire [1:0] _GEN_503 = io_fu_2_valid ? _GEN_473 : _GEN_443; // @[ROB.scala 186:23]
  wire [1:0] _GEN_504 = io_fu_2_valid ? _GEN_474 : _GEN_444; // @[ROB.scala 186:23]
  wire [1:0] _GEN_505 = io_fu_2_valid ? _GEN_475 : _GEN_445; // @[ROB.scala 186:23]
  wire [1:0] _GEN_506 = io_fu_2_valid ? _GEN_476 : _GEN_446; // @[ROB.scala 186:23]
  wire [31:0] _GEN_507 = io_fu_2_valid ? _GEN_477 : _GEN_447; // @[ROB.scala 186:23]
  wire [31:0] _GEN_508 = io_fu_2_valid ? _GEN_478 : _GEN_448; // @[ROB.scala 186:23]
  wire [31:0] _GEN_509 = io_fu_2_valid ? _GEN_479 : _GEN_449; // @[ROB.scala 186:23]
  wire [31:0] _GEN_510 = io_fu_2_valid ? _GEN_480 : _GEN_450; // @[ROB.scala 186:23]
  wire [31:0] _GEN_511 = io_fu_2_valid ? _GEN_481 : _GEN_451; // @[ROB.scala 186:23]
  wire  _GEN_512 = io_fu_2_valid ? _GEN_482 : _GEN_452; // @[ROB.scala 186:23]
  wire  _GEN_513 = io_fu_2_valid ? _GEN_483 : _GEN_453; // @[ROB.scala 186:23]
  wire  _GEN_514 = io_fu_2_valid ? _GEN_484 : _GEN_454; // @[ROB.scala 186:23]
  wire  _GEN_515 = io_fu_2_valid ? _GEN_485 : _GEN_455; // @[ROB.scala 186:23]
  wire  _GEN_516 = io_fu_2_valid ? _GEN_486 : _GEN_456; // @[ROB.scala 186:23]
  wire [31:0] _GEN_517 = io_fu_2_valid ? _GEN_487 : _GEN_457; // @[ROB.scala 186:23]
  wire [31:0] _GEN_518 = io_fu_2_valid ? _GEN_488 : _GEN_458; // @[ROB.scala 186:23]
  wire [31:0] _GEN_519 = io_fu_2_valid ? _GEN_489 : _GEN_459; // @[ROB.scala 186:23]
  wire [31:0] _GEN_520 = io_fu_2_valid ? _GEN_490 : _GEN_460; // @[ROB.scala 186:23]
  wire [31:0] _GEN_521 = io_fu_2_valid ? _GEN_491 : _GEN_461; // @[ROB.scala 186:23]
  wire  _GEN_522 = io_fu_2_valid ? _GEN_492 : _GEN_462; // @[ROB.scala 186:23]
  wire  _GEN_523 = io_fu_2_valid ? _GEN_493 : _GEN_463; // @[ROB.scala 186:23]
  wire  _GEN_524 = io_fu_2_valid ? _GEN_494 : _GEN_464; // @[ROB.scala 186:23]
  wire  _GEN_525 = io_fu_2_valid ? _GEN_495 : _GEN_465; // @[ROB.scala 186:23]
  wire  _GEN_526 = io_fu_2_valid ? _GEN_496 : _GEN_466; // @[ROB.scala 186:23]
  wire [2:0] _T_53 = io_fu_3_bits_id - 3'h1; // @[ROB.scala 187:31]
  wire [1:0] _GEN_532 = 3'h0 == _T_53 ? 2'h2 : _GEN_502; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_533 = 3'h1 == _T_53 ? 2'h2 : _GEN_503; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_534 = 3'h2 == _T_53 ? 2'h2 : _GEN_504; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_535 = 3'h3 == _T_53 ? 2'h2 : _GEN_505; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_536 = 3'h4 == _T_53 ? 2'h2 : _GEN_506; // @[ROB.scala 188:{44,44}]
  wire [1:0] _GEN_562 = io_fu_3_valid ? _GEN_532 : _GEN_502; // @[ROB.scala 186:23]
  wire [1:0] _GEN_563 = io_fu_3_valid ? _GEN_533 : _GEN_503; // @[ROB.scala 186:23]
  wire [1:0] _GEN_564 = io_fu_3_valid ? _GEN_534 : _GEN_504; // @[ROB.scala 186:23]
  wire [1:0] _GEN_565 = io_fu_3_valid ? _GEN_535 : _GEN_505; // @[ROB.scala 186:23]
  wire [1:0] _GEN_566 = io_fu_3_valid ? _GEN_536 : _GEN_506; // @[ROB.scala 186:23]
  wire [2:0] _T_65 = io_rs_0_bits_id - 3'h1; // @[ROB.scala 206:31]
  wire [1:0] _GEN_587 = 3'h0 == _T_65 ? 2'h1 : _GEN_562; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_588 = 3'h1 == _T_65 ? 2'h1 : _GEN_563; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_589 = 3'h2 == _T_65 ? 2'h1 : _GEN_564; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_590 = 3'h3 == _T_65 ? 2'h1 : _GEN_565; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_591 = 3'h4 == _T_65 ? 2'h1 : _GEN_566; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_592 = io_rs_0_valid ? _GEN_587 : _GEN_562; // @[ROB.scala 205:22]
  wire [1:0] _GEN_593 = io_rs_0_valid ? _GEN_588 : _GEN_563; // @[ROB.scala 205:22]
  wire [1:0] _GEN_594 = io_rs_0_valid ? _GEN_589 : _GEN_564; // @[ROB.scala 205:22]
  wire [1:0] _GEN_595 = io_rs_0_valid ? _GEN_590 : _GEN_565; // @[ROB.scala 205:22]
  wire [1:0] _GEN_596 = io_rs_0_valid ? _GEN_591 : _GEN_566; // @[ROB.scala 205:22]
  wire [2:0] _T_67 = io_rs_1_bits_id - 3'h1; // @[ROB.scala 206:31]
  wire [1:0] _GEN_597 = 3'h0 == _T_67 ? 2'h1 : _GEN_592; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_598 = 3'h1 == _T_67 ? 2'h1 : _GEN_593; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_599 = 3'h2 == _T_67 ? 2'h1 : _GEN_594; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_600 = 3'h3 == _T_67 ? 2'h1 : _GEN_595; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_601 = 3'h4 == _T_67 ? 2'h1 : _GEN_596; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_602 = io_rs_1_valid ? _GEN_597 : _GEN_592; // @[ROB.scala 205:22]
  wire [1:0] _GEN_603 = io_rs_1_valid ? _GEN_598 : _GEN_593; // @[ROB.scala 205:22]
  wire [1:0] _GEN_604 = io_rs_1_valid ? _GEN_599 : _GEN_594; // @[ROB.scala 205:22]
  wire [1:0] _GEN_605 = io_rs_1_valid ? _GEN_600 : _GEN_595; // @[ROB.scala 205:22]
  wire [1:0] _GEN_606 = io_rs_1_valid ? _GEN_601 : _GEN_596; // @[ROB.scala 205:22]
  wire [2:0] _T_69 = io_rs_2_bits_id - 3'h1; // @[ROB.scala 206:31]
  wire [1:0] _GEN_607 = 3'h0 == _T_69 ? 2'h1 : _GEN_602; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_608 = 3'h1 == _T_69 ? 2'h1 : _GEN_603; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_609 = 3'h2 == _T_69 ? 2'h1 : _GEN_604; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_610 = 3'h3 == _T_69 ? 2'h1 : _GEN_605; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_611 = 3'h4 == _T_69 ? 2'h1 : _GEN_606; // @[ROB.scala 206:{44,44}]
  wire [1:0] _GEN_612 = io_rs_2_valid ? _GEN_607 : _GEN_602; // @[ROB.scala 205:22]
  wire [1:0] _GEN_613 = io_rs_2_valid ? _GEN_608 : _GEN_603; // @[ROB.scala 205:22]
  wire [1:0] _GEN_614 = io_rs_2_valid ? _GEN_609 : _GEN_604; // @[ROB.scala 205:22]
  wire [1:0] _GEN_615 = io_rs_2_valid ? _GEN_610 : _GEN_605; // @[ROB.scala 205:22]
  wire [1:0] _GEN_616 = io_rs_2_valid ? _GEN_611 : _GEN_606; // @[ROB.scala 205:22]
  wire [2:0] _T_71 = io_rs_3_bits_id - 3'h1; // @[ROB.scala 206:31]
  assign io_enq_ready = ~full & ~_GEN_4; // @[ROB.scala 134:27]
  assign io_deq_valid = _GEN_9 == 2'h2 & _GEN_14; // @[ROB.scala 135:52]
  assign io_deq_bits_rdWrEn = _GEN_24 != 5'h0; // @[ROB.scala 138:44]
  assign io_deq_bits_rd = 3'h4 == head ? entries_4_rd : _GEN_23; // @[ROB.scala 137:{20,20}]
  assign io_deq_bits_data = 3'h4 == head ? entries_4_data : _GEN_18; // @[ROB.scala 136:{22,22}]
  assign io_deq_bits_id = {{5'd0}, _io_deq_bits_id_T_1}; // @[ROB.scala 145:20]
  assign io_deq_bits_brAddr = 3'h4 == head ? entries_4_brAddr : _GEN_38; // @[ROB.scala 141:{24,24}]
  assign io_deq_bits_brTaken = 3'h4 == head ? entries_4_brTaken : _GEN_43; // @[ROB.scala 142:{25,25}]
  assign io_deq_bits_excpAddr = 3'h4 == head ? entries_4_excpAddr : _GEN_48; // @[ROB.scala 143:{26,26}]
  assign io_deq_bits_excpValid = 3'h4 == head ? entries_4_excpValid : _GEN_53; // @[ROB.scala 144:{27,27}]
  assign io_deq_bits_pc = 3'h4 == head ? entries_4_pc : _GEN_28; // @[ROB.scala 139:{20,20}]
  assign io_deq_bits_inst = 3'h4 == head ? entries_4_inst : _GEN_33; // @[ROB.scala 140:{22,22}]
  assign io_read_0_busy = entries_0_busy; // @[ROB.scala 197:16]
  assign io_read_0_state = entries_0_state; // @[ROB.scala 199:17]
  assign io_read_0_rd = entries_0_rd; // @[ROB.scala 200:14]
  assign io_read_0_data = entries_0_data; // @[ROB.scala 198:16]
  assign io_read_1_busy = entries_1_busy; // @[ROB.scala 197:16]
  assign io_read_1_state = entries_1_state; // @[ROB.scala 199:17]
  assign io_read_1_rd = entries_1_rd; // @[ROB.scala 200:14]
  assign io_read_1_data = entries_1_data; // @[ROB.scala 198:16]
  assign io_read_2_busy = entries_2_busy; // @[ROB.scala 197:16]
  assign io_read_2_state = entries_2_state; // @[ROB.scala 199:17]
  assign io_read_2_rd = entries_2_rd; // @[ROB.scala 200:14]
  assign io_read_2_data = entries_2_data; // @[ROB.scala 198:16]
  assign io_read_3_busy = entries_3_busy; // @[ROB.scala 197:16]
  assign io_read_3_state = entries_3_state; // @[ROB.scala 199:17]
  assign io_read_3_rd = entries_3_rd; // @[ROB.scala 200:14]
  assign io_read_3_data = entries_3_data; // @[ROB.scala 198:16]
  assign io_read_4_busy = entries_4_busy; // @[ROB.scala 197:16]
  assign io_read_4_state = entries_4_state; // @[ROB.scala 199:17]
  assign io_read_4_rd = entries_4_rd; // @[ROB.scala 200:14]
  assign io_read_4_data = entries_4_data; // @[ROB.scala 198:16]
  assign io_id = tail + 3'h1; // @[ROB.scala 133:19]
  assign io_regStatus_0_owner = regResStat_0_owner; // @[ROB.scala 132:18]
  assign io_regStatus_1_owner = regResStat_1_owner; // @[ROB.scala 132:18]
  assign io_regStatus_2_owner = regResStat_2_owner; // @[ROB.scala 132:18]
  assign io_regStatus_3_owner = regResStat_3_owner; // @[ROB.scala 132:18]
  assign io_regStatus_4_owner = regResStat_4_owner; // @[ROB.scala 132:18]
  assign io_regStatus_5_owner = regResStat_5_owner; // @[ROB.scala 132:18]
  assign io_regStatus_6_owner = regResStat_6_owner; // @[ROB.scala 132:18]
  assign io_regStatus_7_owner = regResStat_7_owner; // @[ROB.scala 132:18]
  assign io_regStatus_8_owner = regResStat_8_owner; // @[ROB.scala 132:18]
  assign io_regStatus_9_owner = regResStat_9_owner; // @[ROB.scala 132:18]
  assign io_regStatus_10_owner = regResStat_10_owner; // @[ROB.scala 132:18]
  assign io_regStatus_11_owner = regResStat_11_owner; // @[ROB.scala 132:18]
  assign io_regStatus_12_owner = regResStat_12_owner; // @[ROB.scala 132:18]
  assign io_regStatus_13_owner = regResStat_13_owner; // @[ROB.scala 132:18]
  assign io_regStatus_14_owner = regResStat_14_owner; // @[ROB.scala 132:18]
  assign io_regStatus_15_owner = regResStat_15_owner; // @[ROB.scala 132:18]
  assign io_regStatus_16_owner = regResStat_16_owner; // @[ROB.scala 132:18]
  assign io_regStatus_17_owner = regResStat_17_owner; // @[ROB.scala 132:18]
  assign io_regStatus_18_owner = regResStat_18_owner; // @[ROB.scala 132:18]
  assign io_regStatus_19_owner = regResStat_19_owner; // @[ROB.scala 132:18]
  assign io_regStatus_20_owner = regResStat_20_owner; // @[ROB.scala 132:18]
  assign io_regStatus_21_owner = regResStat_21_owner; // @[ROB.scala 132:18]
  assign io_regStatus_22_owner = regResStat_22_owner; // @[ROB.scala 132:18]
  assign io_regStatus_23_owner = regResStat_23_owner; // @[ROB.scala 132:18]
  assign io_regStatus_24_owner = regResStat_24_owner; // @[ROB.scala 132:18]
  assign io_regStatus_25_owner = regResStat_25_owner; // @[ROB.scala 132:18]
  assign io_regStatus_26_owner = regResStat_26_owner; // @[ROB.scala 132:18]
  assign io_regStatus_27_owner = regResStat_27_owner; // @[ROB.scala 132:18]
  assign io_regStatus_28_owner = regResStat_28_owner; // @[ROB.scala 132:18]
  assign io_regStatus_29_owner = regResStat_29_owner; // @[ROB.scala 132:18]
  assign io_regStatus_30_owner = regResStat_30_owner; // @[ROB.scala 132:18]
  assign io_regStatus_31_owner = regResStat_31_owner; // @[ROB.scala 132:18]
  always @(posedge clock) begin
    if (io_flush) begin // @[ROB.scala 210:21]
      entries_0_busy <= 1'h0; // @[ROB.scala 211:37]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (3'h0 == head) begin // @[ROB.scala 163:28]
        entries_0_busy <= 1'h0; // @[ROB.scala 163:28]
      end else begin
        entries_0_busy <= _GEN_117;
      end
    end else begin
      entries_0_busy <= _GEN_117;
    end
    if (io_rs_3_valid) begin // @[ROB.scala 205:22]
      if (3'h0 == _T_71) begin // @[ROB.scala 206:44]
        entries_0_state <= 2'h1; // @[ROB.scala 206:44]
      end else begin
        entries_0_state <= _GEN_612;
      end
    end else begin
      entries_0_state <= _GEN_612;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h0 == tail) begin // @[ROB.scala 152:26]
        entries_0_rd <= io_enq_bits_rd; // @[ROB.scala 152:26]
      end
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h0 == _T_53) begin // @[ROB.scala 187:43]
        entries_0_data <= io_fu_3_bits_data; // @[ROB.scala 187:43]
      end else begin
        entries_0_data <= _GEN_497;
      end
    end else begin
      entries_0_data <= _GEN_497;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h0 == _T_53) begin // @[ROB.scala 189:45]
        entries_0_brAddr <= 32'h0; // @[ROB.scala 189:45]
      end else begin
        entries_0_brAddr <= _GEN_507;
      end
    end else begin
      entries_0_brAddr <= _GEN_507;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h0 == _T_53) begin // @[ROB.scala 190:46]
        entries_0_brTaken <= 1'h0; // @[ROB.scala 190:46]
      end else begin
        entries_0_brTaken <= _GEN_512;
      end
    end else begin
      entries_0_brTaken <= _GEN_512;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h0 == _T_53) begin // @[ROB.scala 191:47]
        entries_0_excpAddr <= io_fu_3_bits_excpAddr; // @[ROB.scala 191:47]
      end else begin
        entries_0_excpAddr <= _GEN_517;
      end
    end else begin
      entries_0_excpAddr <= _GEN_517;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h0 == _T_53) begin // @[ROB.scala 192:48]
        entries_0_excpValid <= io_fu_3_bits_excpValid; // @[ROB.scala 192:48]
      end else begin
        entries_0_excpValid <= _GEN_522;
      end
    end else begin
      entries_0_excpValid <= _GEN_522;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h0 == tail) begin // @[ROB.scala 153:26]
        entries_0_pc <= io_enq_bits_pc; // @[ROB.scala 153:26]
      end
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h0 == tail) begin // @[ROB.scala 154:28]
        entries_0_inst <= io_enq_bits_inst; // @[ROB.scala 154:28]
      end
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      entries_1_busy <= 1'h0; // @[ROB.scala 211:37]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (3'h1 == head) begin // @[ROB.scala 163:28]
        entries_1_busy <= 1'h0; // @[ROB.scala 163:28]
      end else begin
        entries_1_busy <= _GEN_118;
      end
    end else begin
      entries_1_busy <= _GEN_118;
    end
    if (io_rs_3_valid) begin // @[ROB.scala 205:22]
      if (3'h1 == _T_71) begin // @[ROB.scala 206:44]
        entries_1_state <= 2'h1; // @[ROB.scala 206:44]
      end else begin
        entries_1_state <= _GEN_613;
      end
    end else begin
      entries_1_state <= _GEN_613;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h1 == tail) begin // @[ROB.scala 152:26]
        entries_1_rd <= io_enq_bits_rd; // @[ROB.scala 152:26]
      end
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h1 == _T_53) begin // @[ROB.scala 187:43]
        entries_1_data <= io_fu_3_bits_data; // @[ROB.scala 187:43]
      end else begin
        entries_1_data <= _GEN_498;
      end
    end else begin
      entries_1_data <= _GEN_498;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h1 == _T_53) begin // @[ROB.scala 189:45]
        entries_1_brAddr <= 32'h0; // @[ROB.scala 189:45]
      end else begin
        entries_1_brAddr <= _GEN_508;
      end
    end else begin
      entries_1_brAddr <= _GEN_508;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h1 == _T_53) begin // @[ROB.scala 190:46]
        entries_1_brTaken <= 1'h0; // @[ROB.scala 190:46]
      end else begin
        entries_1_brTaken <= _GEN_513;
      end
    end else begin
      entries_1_brTaken <= _GEN_513;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h1 == _T_53) begin // @[ROB.scala 191:47]
        entries_1_excpAddr <= io_fu_3_bits_excpAddr; // @[ROB.scala 191:47]
      end else begin
        entries_1_excpAddr <= _GEN_518;
      end
    end else begin
      entries_1_excpAddr <= _GEN_518;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h1 == _T_53) begin // @[ROB.scala 192:48]
        entries_1_excpValid <= io_fu_3_bits_excpValid; // @[ROB.scala 192:48]
      end else begin
        entries_1_excpValid <= _GEN_523;
      end
    end else begin
      entries_1_excpValid <= _GEN_523;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h1 == tail) begin // @[ROB.scala 153:26]
        entries_1_pc <= io_enq_bits_pc; // @[ROB.scala 153:26]
      end
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h1 == tail) begin // @[ROB.scala 154:28]
        entries_1_inst <= io_enq_bits_inst; // @[ROB.scala 154:28]
      end
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      entries_2_busy <= 1'h0; // @[ROB.scala 211:37]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (3'h2 == head) begin // @[ROB.scala 163:28]
        entries_2_busy <= 1'h0; // @[ROB.scala 163:28]
      end else begin
        entries_2_busy <= _GEN_119;
      end
    end else begin
      entries_2_busy <= _GEN_119;
    end
    if (io_rs_3_valid) begin // @[ROB.scala 205:22]
      if (3'h2 == _T_71) begin // @[ROB.scala 206:44]
        entries_2_state <= 2'h1; // @[ROB.scala 206:44]
      end else begin
        entries_2_state <= _GEN_614;
      end
    end else begin
      entries_2_state <= _GEN_614;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h2 == tail) begin // @[ROB.scala 152:26]
        entries_2_rd <= io_enq_bits_rd; // @[ROB.scala 152:26]
      end
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h2 == _T_53) begin // @[ROB.scala 187:43]
        entries_2_data <= io_fu_3_bits_data; // @[ROB.scala 187:43]
      end else begin
        entries_2_data <= _GEN_499;
      end
    end else begin
      entries_2_data <= _GEN_499;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h2 == _T_53) begin // @[ROB.scala 189:45]
        entries_2_brAddr <= 32'h0; // @[ROB.scala 189:45]
      end else begin
        entries_2_brAddr <= _GEN_509;
      end
    end else begin
      entries_2_brAddr <= _GEN_509;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h2 == _T_53) begin // @[ROB.scala 190:46]
        entries_2_brTaken <= 1'h0; // @[ROB.scala 190:46]
      end else begin
        entries_2_brTaken <= _GEN_514;
      end
    end else begin
      entries_2_brTaken <= _GEN_514;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h2 == _T_53) begin // @[ROB.scala 191:47]
        entries_2_excpAddr <= io_fu_3_bits_excpAddr; // @[ROB.scala 191:47]
      end else begin
        entries_2_excpAddr <= _GEN_519;
      end
    end else begin
      entries_2_excpAddr <= _GEN_519;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h2 == _T_53) begin // @[ROB.scala 192:48]
        entries_2_excpValid <= io_fu_3_bits_excpValid; // @[ROB.scala 192:48]
      end else begin
        entries_2_excpValid <= _GEN_524;
      end
    end else begin
      entries_2_excpValid <= _GEN_524;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h2 == tail) begin // @[ROB.scala 153:26]
        entries_2_pc <= io_enq_bits_pc; // @[ROB.scala 153:26]
      end
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h2 == tail) begin // @[ROB.scala 154:28]
        entries_2_inst <= io_enq_bits_inst; // @[ROB.scala 154:28]
      end
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      entries_3_busy <= 1'h0; // @[ROB.scala 211:37]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (3'h3 == head) begin // @[ROB.scala 163:28]
        entries_3_busy <= 1'h0; // @[ROB.scala 163:28]
      end else begin
        entries_3_busy <= _GEN_120;
      end
    end else begin
      entries_3_busy <= _GEN_120;
    end
    if (io_rs_3_valid) begin // @[ROB.scala 205:22]
      if (3'h3 == _T_71) begin // @[ROB.scala 206:44]
        entries_3_state <= 2'h1; // @[ROB.scala 206:44]
      end else begin
        entries_3_state <= _GEN_615;
      end
    end else begin
      entries_3_state <= _GEN_615;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h3 == tail) begin // @[ROB.scala 152:26]
        entries_3_rd <= io_enq_bits_rd; // @[ROB.scala 152:26]
      end
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h3 == _T_53) begin // @[ROB.scala 187:43]
        entries_3_data <= io_fu_3_bits_data; // @[ROB.scala 187:43]
      end else begin
        entries_3_data <= _GEN_500;
      end
    end else begin
      entries_3_data <= _GEN_500;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h3 == _T_53) begin // @[ROB.scala 189:45]
        entries_3_brAddr <= 32'h0; // @[ROB.scala 189:45]
      end else begin
        entries_3_brAddr <= _GEN_510;
      end
    end else begin
      entries_3_brAddr <= _GEN_510;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h3 == _T_53) begin // @[ROB.scala 190:46]
        entries_3_brTaken <= 1'h0; // @[ROB.scala 190:46]
      end else begin
        entries_3_brTaken <= _GEN_515;
      end
    end else begin
      entries_3_brTaken <= _GEN_515;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h3 == _T_53) begin // @[ROB.scala 191:47]
        entries_3_excpAddr <= io_fu_3_bits_excpAddr; // @[ROB.scala 191:47]
      end else begin
        entries_3_excpAddr <= _GEN_520;
      end
    end else begin
      entries_3_excpAddr <= _GEN_520;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h3 == _T_53) begin // @[ROB.scala 192:48]
        entries_3_excpValid <= io_fu_3_bits_excpValid; // @[ROB.scala 192:48]
      end else begin
        entries_3_excpValid <= _GEN_525;
      end
    end else begin
      entries_3_excpValid <= _GEN_525;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h3 == tail) begin // @[ROB.scala 153:26]
        entries_3_pc <= io_enq_bits_pc; // @[ROB.scala 153:26]
      end
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h3 == tail) begin // @[ROB.scala 154:28]
        entries_3_inst <= io_enq_bits_inst; // @[ROB.scala 154:28]
      end
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      entries_4_busy <= 1'h0; // @[ROB.scala 211:37]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (3'h4 == head) begin // @[ROB.scala 163:28]
        entries_4_busy <= 1'h0; // @[ROB.scala 163:28]
      end else begin
        entries_4_busy <= _GEN_121;
      end
    end else begin
      entries_4_busy <= _GEN_121;
    end
    if (io_rs_3_valid) begin // @[ROB.scala 205:22]
      if (3'h4 == _T_71) begin // @[ROB.scala 206:44]
        entries_4_state <= 2'h1; // @[ROB.scala 206:44]
      end else begin
        entries_4_state <= _GEN_616;
      end
    end else begin
      entries_4_state <= _GEN_616;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h4 == tail) begin // @[ROB.scala 152:26]
        entries_4_rd <= io_enq_bits_rd; // @[ROB.scala 152:26]
      end
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h4 == _T_53) begin // @[ROB.scala 187:43]
        entries_4_data <= io_fu_3_bits_data; // @[ROB.scala 187:43]
      end else begin
        entries_4_data <= _GEN_501;
      end
    end else begin
      entries_4_data <= _GEN_501;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h4 == _T_53) begin // @[ROB.scala 189:45]
        entries_4_brAddr <= 32'h0; // @[ROB.scala 189:45]
      end else begin
        entries_4_brAddr <= _GEN_511;
      end
    end else begin
      entries_4_brAddr <= _GEN_511;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h4 == _T_53) begin // @[ROB.scala 190:46]
        entries_4_brTaken <= 1'h0; // @[ROB.scala 190:46]
      end else begin
        entries_4_brTaken <= _GEN_516;
      end
    end else begin
      entries_4_brTaken <= _GEN_516;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h4 == _T_53) begin // @[ROB.scala 191:47]
        entries_4_excpAddr <= io_fu_3_bits_excpAddr; // @[ROB.scala 191:47]
      end else begin
        entries_4_excpAddr <= _GEN_521;
      end
    end else begin
      entries_4_excpAddr <= _GEN_521;
    end
    if (io_fu_3_valid) begin // @[ROB.scala 186:23]
      if (3'h4 == _T_53) begin // @[ROB.scala 192:48]
        entries_4_excpValid <= io_fu_3_bits_excpValid; // @[ROB.scala 192:48]
      end else begin
        entries_4_excpValid <= _GEN_526;
      end
    end else begin
      entries_4_excpValid <= _GEN_526;
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h4 == tail) begin // @[ROB.scala 153:26]
        entries_4_pc <= io_enq_bits_pc; // @[ROB.scala 153:26]
      end
    end
    if (_T) begin // @[ROB.scala 148:24]
      if (3'h4 == tail) begin // @[ROB.scala 154:28]
        entries_4_inst <= io_enq_bits_inst; // @[ROB.scala 154:28]
      end
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_0_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h0 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_0_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_0_owner <= _GEN_142;
        end
      end else begin
        regResStat_0_owner <= _GEN_142;
      end
    end else begin
      regResStat_0_owner <= _GEN_142;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_1_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h1 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_1_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_1_owner <= _GEN_143;
        end
      end else begin
        regResStat_1_owner <= _GEN_143;
      end
    end else begin
      regResStat_1_owner <= _GEN_143;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_2_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h2 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_2_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_2_owner <= _GEN_144;
        end
      end else begin
        regResStat_2_owner <= _GEN_144;
      end
    end else begin
      regResStat_2_owner <= _GEN_144;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_3_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h3 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_3_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_3_owner <= _GEN_145;
        end
      end else begin
        regResStat_3_owner <= _GEN_145;
      end
    end else begin
      regResStat_3_owner <= _GEN_145;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_4_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h4 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_4_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_4_owner <= _GEN_146;
        end
      end else begin
        regResStat_4_owner <= _GEN_146;
      end
    end else begin
      regResStat_4_owner <= _GEN_146;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_5_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h5 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_5_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_5_owner <= _GEN_147;
        end
      end else begin
        regResStat_5_owner <= _GEN_147;
      end
    end else begin
      regResStat_5_owner <= _GEN_147;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_6_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h6 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_6_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_6_owner <= _GEN_148;
        end
      end else begin
        regResStat_6_owner <= _GEN_148;
      end
    end else begin
      regResStat_6_owner <= _GEN_148;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_7_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h7 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_7_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_7_owner <= _GEN_149;
        end
      end else begin
        regResStat_7_owner <= _GEN_149;
      end
    end else begin
      regResStat_7_owner <= _GEN_149;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_8_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h8 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_8_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_8_owner <= _GEN_150;
        end
      end else begin
        regResStat_8_owner <= _GEN_150;
      end
    end else begin
      regResStat_8_owner <= _GEN_150;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_9_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h9 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_9_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_9_owner <= _GEN_151;
        end
      end else begin
        regResStat_9_owner <= _GEN_151;
      end
    end else begin
      regResStat_9_owner <= _GEN_151;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_10_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'ha == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_10_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_10_owner <= _GEN_152;
        end
      end else begin
        regResStat_10_owner <= _GEN_152;
      end
    end else begin
      regResStat_10_owner <= _GEN_152;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_11_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'hb == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_11_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_11_owner <= _GEN_153;
        end
      end else begin
        regResStat_11_owner <= _GEN_153;
      end
    end else begin
      regResStat_11_owner <= _GEN_153;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_12_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'hc == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_12_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_12_owner <= _GEN_154;
        end
      end else begin
        regResStat_12_owner <= _GEN_154;
      end
    end else begin
      regResStat_12_owner <= _GEN_154;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_13_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'hd == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_13_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_13_owner <= _GEN_155;
        end
      end else begin
        regResStat_13_owner <= _GEN_155;
      end
    end else begin
      regResStat_13_owner <= _GEN_155;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_14_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'he == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_14_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_14_owner <= _GEN_156;
        end
      end else begin
        regResStat_14_owner <= _GEN_156;
      end
    end else begin
      regResStat_14_owner <= _GEN_156;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_15_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'hf == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_15_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_15_owner <= _GEN_157;
        end
      end else begin
        regResStat_15_owner <= _GEN_157;
      end
    end else begin
      regResStat_15_owner <= _GEN_157;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_16_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h10 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_16_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_16_owner <= _GEN_158;
        end
      end else begin
        regResStat_16_owner <= _GEN_158;
      end
    end else begin
      regResStat_16_owner <= _GEN_158;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_17_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h11 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_17_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_17_owner <= _GEN_159;
        end
      end else begin
        regResStat_17_owner <= _GEN_159;
      end
    end else begin
      regResStat_17_owner <= _GEN_159;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_18_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h12 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_18_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_18_owner <= _GEN_160;
        end
      end else begin
        regResStat_18_owner <= _GEN_160;
      end
    end else begin
      regResStat_18_owner <= _GEN_160;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_19_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h13 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_19_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_19_owner <= _GEN_161;
        end
      end else begin
        regResStat_19_owner <= _GEN_161;
      end
    end else begin
      regResStat_19_owner <= _GEN_161;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_20_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h14 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_20_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_20_owner <= _GEN_162;
        end
      end else begin
        regResStat_20_owner <= _GEN_162;
      end
    end else begin
      regResStat_20_owner <= _GEN_162;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_21_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h15 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_21_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_21_owner <= _GEN_163;
        end
      end else begin
        regResStat_21_owner <= _GEN_163;
      end
    end else begin
      regResStat_21_owner <= _GEN_163;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_22_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h16 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_22_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_22_owner <= _GEN_164;
        end
      end else begin
        regResStat_22_owner <= _GEN_164;
      end
    end else begin
      regResStat_22_owner <= _GEN_164;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_23_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h17 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_23_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_23_owner <= _GEN_165;
        end
      end else begin
        regResStat_23_owner <= _GEN_165;
      end
    end else begin
      regResStat_23_owner <= _GEN_165;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_24_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h18 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_24_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_24_owner <= _GEN_166;
        end
      end else begin
        regResStat_24_owner <= _GEN_166;
      end
    end else begin
      regResStat_24_owner <= _GEN_166;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_25_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h19 == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_25_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_25_owner <= _GEN_167;
        end
      end else begin
        regResStat_25_owner <= _GEN_167;
      end
    end else begin
      regResStat_25_owner <= _GEN_167;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_26_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h1a == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_26_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_26_owner <= _GEN_168;
        end
      end else begin
        regResStat_26_owner <= _GEN_168;
      end
    end else begin
      regResStat_26_owner <= _GEN_168;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_27_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h1b == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_27_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_27_owner <= _GEN_169;
        end
      end else begin
        regResStat_27_owner <= _GEN_169;
      end
    end else begin
      regResStat_27_owner <= _GEN_169;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_28_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h1c == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_28_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_28_owner <= _GEN_170;
        end
      end else begin
        regResStat_28_owner <= _GEN_170;
      end
    end else begin
      regResStat_28_owner <= _GEN_170;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_29_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h1d == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_29_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_29_owner <= _GEN_171;
        end
      end else begin
        regResStat_29_owner <= _GEN_171;
      end
    end else begin
      regResStat_29_owner <= _GEN_171;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_30_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h1e == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_30_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_30_owner <= _GEN_172;
        end
      end else begin
        regResStat_30_owner <= _GEN_172;
      end
    end else begin
      regResStat_30_owner <= _GEN_172;
    end
    if (io_flush) begin // @[ROB.scala 210:21]
      regResStat_31_owner <= 8'h0; // @[ROB.scala 212:41]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (_GEN_226 == _GEN_672 & ~(_T & io_enq_bits_rd == _GEN_24)) begin // @[ROB.scala 169:111]
        if (5'h1f == _GEN_24) begin // @[ROB.scala 170:42]
          regResStat_31_owner <= 8'h0; // @[ROB.scala 170:42]
        end else begin
          regResStat_31_owner <= _GEN_173;
        end
      end else begin
        regResStat_31_owner <= _GEN_173;
      end
    end else begin
      regResStat_31_owner <= _GEN_173;
    end
    if (reset) begin // @[ROB.scala 121:23]
      head <= 3'h0; // @[ROB.scala 121:23]
    end else if (io_flush) begin // @[ROB.scala 210:21]
      head <= 3'h0; // @[ROB.scala 213:14]
    end else if (io_deq_valid) begin // @[ROB.scala 162:24]
      if (head == 3'h4) begin // @[ROB.scala 173:20]
        head <= 3'h0;
      end else begin
        head <= _io_deq_bits_id_T_1;
      end
    end
    if (reset) begin // @[ROB.scala 122:23]
      tail <= 3'h0; // @[ROB.scala 122:23]
    end else if (io_flush) begin // @[ROB.scala 210:21]
      tail <= 3'h0; // @[ROB.scala 214:14]
    end else if (_T) begin // @[ROB.scala 148:24]
      if (tail == 3'h4) begin // @[ROB.scala 159:20]
        tail <= 3'h0;
      end else begin
        tail <= _io_id_T_1;
      end
    end
    if (reset) begin // @[ROB.scala 124:24]
      count <= 3'h0; // @[ROB.scala 124:24]
    end else if (io_flush) begin // @[ROB.scala 210:21]
      count <= 3'h0; // @[ROB.scala 215:15]
    end else if (~(io_deq_valid & _T)) begin // @[ROB.scala 176:43]
      if (io_deq_valid) begin // @[ROB.scala 180:27]
        count <= _count_T_3; // @[ROB.scala 181:19]
      end else begin
        count <= _GEN_344;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  entries_0_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  entries_0_state = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  entries_0_rd = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  entries_0_data = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  entries_0_brAddr = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  entries_0_brTaken = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  entries_0_excpAddr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  entries_0_excpValid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  entries_0_pc = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  entries_0_inst = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  entries_1_busy = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  entries_1_state = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  entries_1_rd = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  entries_1_data = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  entries_1_brAddr = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  entries_1_brTaken = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  entries_1_excpAddr = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  entries_1_excpValid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  entries_1_pc = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  entries_1_inst = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  entries_2_busy = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  entries_2_state = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  entries_2_rd = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  entries_2_data = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  entries_2_brAddr = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  entries_2_brTaken = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  entries_2_excpAddr = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  entries_2_excpValid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  entries_2_pc = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  entries_2_inst = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  entries_3_busy = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  entries_3_state = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  entries_3_rd = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  entries_3_data = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  entries_3_brAddr = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  entries_3_brTaken = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  entries_3_excpAddr = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  entries_3_excpValid = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  entries_3_pc = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  entries_3_inst = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  entries_4_busy = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  entries_4_state = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  entries_4_rd = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  entries_4_data = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  entries_4_brAddr = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  entries_4_brTaken = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  entries_4_excpAddr = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  entries_4_excpValid = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  entries_4_pc = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  entries_4_inst = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  regResStat_0_owner = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  regResStat_1_owner = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  regResStat_2_owner = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  regResStat_3_owner = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  regResStat_4_owner = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  regResStat_5_owner = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  regResStat_6_owner = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  regResStat_7_owner = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  regResStat_8_owner = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  regResStat_9_owner = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  regResStat_10_owner = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  regResStat_11_owner = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  regResStat_12_owner = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  regResStat_13_owner = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  regResStat_14_owner = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  regResStat_15_owner = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  regResStat_16_owner = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  regResStat_17_owner = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  regResStat_18_owner = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  regResStat_19_owner = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  regResStat_20_owner = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  regResStat_21_owner = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  regResStat_22_owner = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  regResStat_23_owner = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  regResStat_24_owner = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  regResStat_25_owner = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  regResStat_26_owner = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  regResStat_27_owner = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  regResStat_28_owner = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  regResStat_29_owner = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  regResStat_30_owner = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  regResStat_31_owner = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  head = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  tail = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  count = _RAND_84[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ImmGen(
  input  [31:0] io_inst,
  input  [2:0]  io_immSrc,
  input         io_immSign,
  output [31:0] io_imm
);
  wire [31:0] immI = {{20'd0}, io_inst[31:20]}; // @[util.scala 62:36]
  wire [11:0] _immS_T_2 = {io_inst[31:25],io_inst[11:7]}; // @[Cat.scala 33:92]
  wire [31:0] immS = {{20'd0}, _immS_T_2}; // @[util.scala 62:36]
  wire [12:0] _immB_T_4 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] immB = {{19'd0}, _immB_T_4}; // @[util.scala 62:36]
  wire [31:0] immU = {io_inst[31:12], 12'h0}; // @[ImmGen.scala 26:36]
  wire [20:0] _immJ_T_4 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] immJ = {{11'd0}, _immJ_T_4}; // @[util.scala 62:36]
  wire [11:0] _immI_S_T_1 = io_inst[31:20]; // @[util.scala 51:20]
  wire  immI_S_signBit = _immI_S_T_1[11]; // @[util.scala 42:27]
  wire [9:0] immI_S_out_lo = {immI_S_signBit,immI_S_signBit,immI_S_signBit,immI_S_signBit,immI_S_signBit,immI_S_signBit,
    immI_S_signBit,immI_S_signBit,immI_S_signBit,immI_S_signBit}; // @[Cat.scala 33:92]
  wire [11:0] _immI_S_out_T_1 = io_inst[31:20]; // @[util.scala 46:75]
  wire [31:0] immI_S = {immI_S_out_lo,immI_S_out_lo,_immI_S_out_T_1}; // @[Cat.scala 33:92]
  wire [11:0] _immS_S_T_3 = {io_inst[31:25],io_inst[11:7]}; // @[util.scala 51:20]
  wire  immS_S_signBit = _immS_S_T_3[11]; // @[util.scala 42:27]
  wire [9:0] immS_S_out_lo = {immS_S_signBit,immS_S_signBit,immS_S_signBit,immS_S_signBit,immS_S_signBit,immS_S_signBit,
    immS_S_signBit,immS_S_signBit,immS_S_signBit,immS_S_signBit}; // @[Cat.scala 33:92]
  wire [11:0] _immS_S_out_T_1 = {io_inst[31:25],io_inst[11:7]}; // @[util.scala 46:75]
  wire [31:0] immS_S = {immS_S_out_lo,immS_S_out_lo,_immS_S_out_T_1}; // @[Cat.scala 33:92]
  wire [12:0] _immB_S_T_5 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[util.scala 51:20]
  wire  immB_S_signBit = _immB_S_T_5[12]; // @[util.scala 42:27]
  wire [9:0] immB_S_out_hi = {immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,
    immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit}; // @[Cat.scala 33:92]
  wire [18:0] _immB_S_out_T = {immB_S_out_hi,immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,
    immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit}; // @[Cat.scala 33:92]
  wire [12:0] _immB_S_out_T_1 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[util.scala 46:75]
  wire [31:0] immB_S = {_immB_S_out_T,_immB_S_out_T_1}; // @[Cat.scala 33:92]
  wire [31:0] immU_S = {io_inst[31:12], 12'h0}; // @[util.scala 44:18]
  wire [20:0] _immJ_S_T_5 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[util.scala 51:20]
  wire  immJ_S_signBit = _immJ_S_T_5[20]; // @[util.scala 42:27]
  wire [4:0] immJ_S_out_lo = {immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit}; // @[Cat.scala 33:92]
  wire [20:0] _immJ_S_out_T_1 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[util.scala 46:75]
  wire [31:0] immJ_S = {immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,
    immJ_S_out_lo,_immJ_S_out_T_1}; // @[Cat.scala 33:92]
  wire [31:0] _out_T_3 = 3'h1 == io_immSrc ? immS_S : immI_S; // @[Mux.scala 81:58]
  wire [31:0] _out_T_5 = 3'h2 == io_immSrc ? immB_S : _out_T_3; // @[Mux.scala 81:58]
  wire [31:0] _out_T_7 = 3'h3 == io_immSrc ? immU_S : _out_T_5; // @[Mux.scala 81:58]
  wire [31:0] _out_T_9 = 3'h4 == io_immSrc ? immJ_S : _out_T_7; // @[Mux.scala 81:58]
  wire [31:0] _out_T_13 = 3'h1 == io_immSrc ? immS : immI; // @[Mux.scala 81:58]
  wire [31:0] _out_T_15 = 3'h2 == io_immSrc ? immB : _out_T_13; // @[Mux.scala 81:58]
  wire [31:0] _out_T_17 = 3'h3 == io_immSrc ? immU : _out_T_15; // @[Mux.scala 81:58]
  wire [31:0] _out_T_19 = 3'h4 == io_immSrc ? immJ : _out_T_17; // @[Mux.scala 81:58]
  wire [31:0] _GEN_0 = io_immSign ? _out_T_9 : _out_T_19; // @[ImmGen.scala 37:19 38:13 46:13]
  wire [31:0] out_out = {{27'd0}, io_inst[19:15]}; // @[util.scala 62:36]
  assign io_imm = io_immSrc == 3'h5 ? out_out : _GEN_0; // @[ImmGen.scala 55:30 56:13]
endmodule
module ALU_1(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  input  [4:0]  io_opSel,
  output [31:0] io_out
);
  wire [31:0] _sum_T_2 = 32'h0 - io_in2; // @[ALU.scala 28:41]
  wire [31:0] _sum_T_3 = io_opSel[0] ? _sum_T_2 : io_in2; // @[ALU.scala 28:27]
  wire [31:0] sum = io_in1 + _sum_T_3; // @[ALU.scala 28:22]
  wire [4:0] shamt = io_in2[4:0]; // @[ALU.scala 31:23]
  wire [31:0] _shiftr_T_1 = io_in1 >> shamt; // @[ALU.scala 33:32]
  wire [31:0] _shiftr_T_4 = $signed(io_in1) >>> shamt; // @[ALU.scala 34:49]
  wire [31:0] shiftr = io_opSel[1] ? _shiftr_T_1 : _shiftr_T_4; // @[ALU.scala 32:21]
  wire [62:0] _GEN_5 = {{31'd0}, io_in1}; // @[ALU.scala 36:25]
  wire [62:0] shiftl = _GEN_5 << shamt; // @[ALU.scala 36:25]
  wire [31:0] _shout_T_3 = io_opSel == 5'hb | io_opSel == 5'hc ? shiftr : 32'h0; // @[ALU.scala 37:20]
  wire [62:0] _shout_T_5 = io_opSel == 5'ha ? shiftl : 63'h0; // @[ALU.scala 38:20]
  wire [62:0] _GEN_2 = {{31'd0}, _shout_T_3}; // @[ALU.scala 37:80]
  wire [62:0] shout = _GEN_2 | _shout_T_5; // @[ALU.scala 37:80]
  wire [31:0] _logic_T = io_in1 & io_in2; // @[ALU.scala 42:40]
  wire [31:0] _logic_T_1 = io_in1 | io_in2; // @[ALU.scala 43:40]
  wire [31:0] _logic_T_2 = io_in1 ^ io_in2; // @[ALU.scala 44:40]
  wire [31:0] _logic_T_4 = 5'h2 == io_opSel ? _logic_T : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _logic_T_6 = 5'h3 == io_opSel ? _logic_T_1 : _logic_T_4; // @[Mux.scala 81:58]
  wire [31:0] logic_ = 5'h4 == io_opSel ? _logic_T_2 : _logic_T_6; // @[Mux.scala 81:58]
  wire  _cmp_T_2 = $signed(io_in1) < $signed(io_in2); // @[ALU.scala 49:48]
  wire  _cmp_T_3 = io_in1 < io_in2; // @[ALU.scala 50:41]
  wire  _cmp_T_4 = io_in1 == io_in2; // @[ALU.scala 51:41]
  wire  _cmp_T_5 = io_in1 != io_in2; // @[ALU.scala 52:41]
  wire  _cmp_T_8 = $signed(io_in1) >= $signed(io_in2); // @[ALU.scala 53:48]
  wire  _cmp_T_9 = io_in1 >= io_in2; // @[ALU.scala 54:42]
  wire  _cmp_T_13 = 5'h9 == io_opSel ? _cmp_T_3 : 5'h8 == io_opSel & _cmp_T_2; // @[Mux.scala 81:58]
  wire  _cmp_T_15 = 5'h5 == io_opSel ? _cmp_T_4 : _cmp_T_13; // @[Mux.scala 81:58]
  wire  _cmp_T_17 = 5'h6 == io_opSel ? _cmp_T_5 : _cmp_T_15; // @[Mux.scala 81:58]
  wire  _cmp_T_19 = 5'h7 == io_opSel ? _cmp_T_8 : _cmp_T_17; // @[Mux.scala 81:58]
  wire  cmp = 5'hf == io_opSel ? _cmp_T_9 : _cmp_T_19; // @[Mux.scala 81:58]
  wire [62:0] _GEN_3 = {{31'd0}, logic_}; // @[ALU.scala 63:68]
  wire [62:0] _io_out_T_3 = _GEN_3 | shout; // @[ALU.scala 63:68]
  wire [62:0] _GEN_4 = {{62'd0}, cmp}; // @[ALU.scala 63:76]
  wire [62:0] _io_out_T_4 = _io_out_T_3 | _GEN_4; // @[ALU.scala 63:76]
  wire [62:0] _io_out_T_5 = io_opSel == 5'h0 | io_opSel == 5'h1 ? {{31'd0}, sum} : _io_out_T_4; // @[ALU.scala 63:22]
  wire [62:0] _GEN_0 = io_opSel == 5'he ? {{31'd0}, io_in2} : _io_out_T_5; // @[ALU.scala 60:33 61:16 63:16]
  wire [62:0] _GEN_1 = io_opSel == 5'hd ? {{31'd0}, io_in1} : _GEN_0; // @[ALU.scala 58:27 59:16]
  assign io_out = _GEN_1[31:0];
endmodule
module ALUStage_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [3:0]  io_in_bits_opr1,
  input  [3:0]  io_in_bits_opr2,
  input  [4:0]  io_in_bits_aluOp,
  input  [2:0]  io_in_bits_immSrc,
  input         io_in_bits_immSign,
  input  [31:0] io_in_bits_rs1Val,
  input  [31:0] io_in_bits_rs2Val,
  input  [31:0] io_in_bits_inst,
  input  [31:0] io_in_bits_pc,
  input  [7:0]  io_in_bits_id,
  output        io_out_valid,
  output [31:0] io_out_bits_data,
  output [7:0]  io_out_bits_id,
  output [4:0]  io_out_bits_rd,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] immGen_io_inst; // @[ALU.scala 230:24]
  wire [2:0] immGen_io_immSrc; // @[ALU.scala 230:24]
  wire  immGen_io_immSign; // @[ALU.scala 230:24]
  wire [31:0] immGen_io_imm; // @[ALU.scala 230:24]
  wire [31:0] alu_io_in1; // @[ALU.scala 258:21]
  wire [31:0] alu_io_in2; // @[ALU.scala 258:21]
  wire [4:0] alu_io_opSel; // @[ALU.scala 258:21]
  wire [31:0] alu_io_out; // @[ALU.scala 258:21]
  reg  s0_full; // @[ALU.scala 221:26]
  wire  s0_ready = ~s0_full; // @[ALU.scala 224:17]
  wire  s0_latch = io_in_valid & s0_ready; // @[ALU.scala 220:32]
  reg  s1_full; // @[ALU.scala 247:26]
  wire  s1_ready = ~s1_full | io_out_valid; // @[ALU.scala 253:26]
  wire  s0_fire = s0_full & s1_ready; // @[ALU.scala 222:28]
  reg [3:0] s0_info_opr1; // @[Reg.scala 19:16]
  reg [3:0] s0_info_opr2; // @[Reg.scala 19:16]
  reg [4:0] s0_info_aluOp; // @[Reg.scala 19:16]
  reg [2:0] s0_info_immSrc; // @[Reg.scala 19:16]
  reg  s0_info_immSign; // @[Reg.scala 19:16]
  reg [31:0] s0_info_rs1Val; // @[Reg.scala 19:16]
  reg [31:0] s0_info_rs2Val; // @[Reg.scala 19:16]
  reg [31:0] s0_info_inst; // @[Reg.scala 19:16]
  reg [31:0] s0_info_pc; // @[Reg.scala 19:16]
  reg [7:0] s0_info_id; // @[Reg.scala 19:16]
  wire  _GEN_10 = s0_fire & s0_full ? 1'h0 : s0_full; // @[ALU.scala 221:26 227:{35,45}]
  wire  _GEN_11 = s0_latch | _GEN_10; // @[ALU.scala 226:{20,30}]
  reg [4:0] s1_rd; // @[Reg.scala 19:16]
  reg [4:0] s1_aluOp; // @[Reg.scala 19:16]
  reg [31:0] s1_aluInVec_0; // @[Reg.scala 19:16]
  reg [31:0] s1_aluInVec_1; // @[Reg.scala 19:16]
  reg [7:0] s1_id; // @[Reg.scala 19:16]
  wire  _GEN_17 = io_out_valid & s1_full ? 1'h0 : s1_full; // @[ALU.scala 247:26 256:{35,45}]
  wire  _GEN_18 = s0_fire | _GEN_17; // @[ALU.scala 255:{20,30}]
  ImmGen immGen ( // @[ALU.scala 230:24]
    .io_inst(immGen_io_inst),
    .io_immSrc(immGen_io_immSrc),
    .io_immSign(immGen_io_immSign),
    .io_imm(immGen_io_imm)
  );
  ALU_1 alu ( // @[ALU.scala 258:21]
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_opSel(alu_io_opSel),
    .io_out(alu_io_out)
  );
  assign io_in_ready = ~s0_full; // @[ALU.scala 224:17]
  assign io_out_valid = s1_full; // @[ALU.scala 266:18]
  assign io_out_bits_data = alu_io_out; // @[ALU.scala 263:22]
  assign io_out_bits_id = s1_id; // @[ALU.scala 264:20]
  assign io_out_bits_rd = s1_rd; // @[ALU.scala 265:20]
  assign immGen_io_inst = s0_info_inst; // @[ALU.scala 234:20]
  assign immGen_io_immSrc = s0_info_immSrc; // @[ALU.scala 232:22]
  assign immGen_io_immSign = s0_info_immSign; // @[ALU.scala 233:23]
  assign alu_io_in1 = s1_aluInVec_0; // @[ALU.scala 259:16]
  assign alu_io_in2 = s1_aluInVec_1; // @[ALU.scala 260:16]
  assign alu_io_opSel = s1_aluOp; // @[ALU.scala 261:18]
  always @(posedge clock) begin
    if (reset) begin // @[ALU.scala 221:26]
      s0_full <= 1'h0; // @[ALU.scala 221:26]
    end else if (io_flush) begin // @[ALU.scala 270:20]
      s0_full <= 1'h0; // @[ALU.scala 271:17]
    end else begin
      s0_full <= _GEN_11;
    end
    if (reset) begin // @[ALU.scala 247:26]
      s1_full <= 1'h0; // @[ALU.scala 247:26]
    end else if (io_flush) begin // @[ALU.scala 270:20]
      s1_full <= 1'h0; // @[ALU.scala 272:17]
    end else begin
      s1_full <= _GEN_18;
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_opr1 <= io_in_bits_opr1; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_opr2 <= io_in_bits_opr2; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_aluOp <= io_in_bits_aluOp; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_immSrc <= io_in_bits_immSrc; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_immSign <= io_in_bits_immSign; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_rs1Val <= io_in_bits_rs1Val; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_rs2Val <= io_in_bits_rs2Val; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_inst <= io_in_bits_inst; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_pc <= io_in_bits_pc; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_id <= io_in_bits_id; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rd <= s0_info_inst[11:7]; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_aluOp <= s0_info_aluOp; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      if (s0_info_opr1 == 4'h0) begin // @[ALU.scala 237:26]
        s1_aluInVec_0 <= 32'h0;
      end else if (s0_info_opr1 == 4'h7) begin // @[ALU.scala 237:62]
        s1_aluInVec_0 <= s0_info_pc;
      end else begin
        s1_aluInVec_0 <= s0_info_rs1Val;
      end
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      if (s0_info_opr2 == 4'h0) begin // @[ALU.scala 238:26]
        s1_aluInVec_1 <= 32'h0;
      end else if (s0_info_opr2 == 4'h3) begin // @[ALU.scala 238:62]
        s1_aluInVec_1 <= immGen_io_imm;
      end else begin
        s1_aluInVec_1 <= s0_info_rs2Val;
      end
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_id <= s0_info_id; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s1_full = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s0_info_opr1 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  s0_info_opr2 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  s0_info_aluOp = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  s0_info_immSrc = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  s0_info_immSign = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s0_info_rs1Val = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  s0_info_rs2Val = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  s0_info_inst = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  s0_info_pc = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  s0_info_id = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  s1_rd = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  s1_aluOp = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  s1_aluInVec_0 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  s1_aluInVec_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  s1_id = _RAND_16[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReservationStation(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [7:0]  io_enq_bits_op,
  input  [3:0]  io_enq_bits_opr1,
  input  [3:0]  io_enq_bits_opr2,
  input  [4:0]  io_enq_bits_rs1,
  input  [4:0]  io_enq_bits_rs2,
  input  [7:0]  io_enq_bits_ROBId,
  input  [7:0]  io_enq_bits_rs1ROBId,
  input  [7:0]  io_enq_bits_rs2ROBId,
  input  [2:0]  io_enq_bits_immSrc,
  input         io_enq_bits_immSign,
  input  [3:0]  io_enq_bits_excpType,
  input  [31:0] io_enq_bits_pc,
  input  [31:0] io_enq_bits_inst,
  input         io_deq_ready,
  output        io_deq_valid,
  output [7:0]  io_deq_bits_op,
  output [7:0]  io_deq_bits_ROBId,
  output [3:0]  io_deq_bits_opr1,
  output [3:0]  io_deq_bits_opr2,
  output [31:0] io_deq_bits_rs1Val,
  output [31:0] io_deq_bits_rs2Val,
  output [2:0]  io_deq_bits_immSrc,
  output        io_deq_bits_immSign,
  output [3:0]  io_deq_bits_excpType,
  output [31:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_inst,
  output        io_robOut_valid,
  output [2:0]  io_robOut_bits_id,
  input         io_robRead_0_busy,
  input  [1:0]  io_robRead_0_state,
  input  [4:0]  io_robRead_0_rd,
  input  [31:0] io_robRead_0_data,
  input         io_robRead_1_busy,
  input  [1:0]  io_robRead_1_state,
  input  [4:0]  io_robRead_1_rd,
  input  [31:0] io_robRead_1_data,
  input         io_robRead_2_busy,
  input  [1:0]  io_robRead_2_state,
  input  [4:0]  io_robRead_2_rd,
  input  [31:0] io_robRead_2_data,
  input         io_robRead_3_busy,
  input  [1:0]  io_robRead_3_state,
  input  [4:0]  io_robRead_3_rd,
  input  [31:0] io_robRead_3_data,
  input         io_robRead_4_busy,
  input  [1:0]  io_robRead_4_state,
  input  [4:0]  io_robRead_4_rd,
  input  [31:0] io_robRead_4_data,
  input  [7:0]  io_regStatus_0_owner,
  input  [7:0]  io_regStatus_1_owner,
  input  [7:0]  io_regStatus_2_owner,
  input  [7:0]  io_regStatus_3_owner,
  input  [7:0]  io_regStatus_4_owner,
  input  [7:0]  io_regStatus_5_owner,
  input  [7:0]  io_regStatus_6_owner,
  input  [7:0]  io_regStatus_7_owner,
  input  [7:0]  io_regStatus_8_owner,
  input  [7:0]  io_regStatus_9_owner,
  input  [7:0]  io_regStatus_10_owner,
  input  [7:0]  io_regStatus_11_owner,
  input  [7:0]  io_regStatus_12_owner,
  input  [7:0]  io_regStatus_13_owner,
  input  [7:0]  io_regStatus_14_owner,
  input  [7:0]  io_regStatus_15_owner,
  input  [7:0]  io_regStatus_16_owner,
  input  [7:0]  io_regStatus_17_owner,
  input  [7:0]  io_regStatus_18_owner,
  input  [7:0]  io_regStatus_19_owner,
  input  [7:0]  io_regStatus_20_owner,
  input  [7:0]  io_regStatus_21_owner,
  input  [7:0]  io_regStatus_22_owner,
  input  [7:0]  io_regStatus_23_owner,
  input  [7:0]  io_regStatus_24_owner,
  input  [7:0]  io_regStatus_25_owner,
  input  [7:0]  io_regStatus_26_owner,
  input  [7:0]  io_regStatus_27_owner,
  input  [7:0]  io_regStatus_28_owner,
  input  [7:0]  io_regStatus_29_owner,
  input  [7:0]  io_regStatus_30_owner,
  input  [7:0]  io_regStatus_31_owner,
  input         io_cdb_0_valid,
  input  [31:0] io_cdb_0_bits_data,
  input  [7:0]  io_cdb_0_bits_id,
  input  [4:0]  io_cdb_0_bits_rd,
  input         io_cdb_1_valid,
  input  [31:0] io_cdb_1_bits_data,
  input  [7:0]  io_cdb_1_bits_id,
  input  [4:0]  io_cdb_1_bits_rd,
  input         io_cdb_2_valid,
  input  [31:0] io_cdb_2_bits_data,
  input  [7:0]  io_cdb_2_bits_id,
  input  [4:0]  io_cdb_2_bits_rd,
  input         io_cdb_3_valid,
  input  [31:0] io_cdb_3_bits_data,
  input  [7:0]  io_cdb_3_bits_id,
  input  [4:0]  io_cdb_3_bits_rd,
  output [4:0]  io_rf_0_addr,
  input  [31:0] io_rf_0_data,
  output [4:0]  io_rf_1_addr,
  input  [31:0] io_rf_1_data,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
`endif // RANDOMIZE_REG_INIT
  reg  entries_0_busy; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_0_op; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_0_ROBId; // @[ReservationStation.scala 85:22]
  reg [3:0] entries_0_opr1; // @[ReservationStation.scala 85:22]
  reg [3:0] entries_0_opr2; // @[ReservationStation.scala 85:22]
  reg [4:0] entries_0_rs1; // @[ReservationStation.scala 85:22]
  reg [4:0] entries_0_rs2; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_0_rs1Val; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_0_rs2Val; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_0_rs1ROBId; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_0_rs2ROBId; // @[ReservationStation.scala 85:22]
  reg [2:0] entries_0_immSrc; // @[ReservationStation.scala 85:22]
  reg  entries_0_immSign; // @[ReservationStation.scala 85:22]
  reg [3:0] entries_0_excpType; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_0_pc; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_0_inst; // @[ReservationStation.scala 85:22]
  reg  entries_1_busy; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_1_op; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_1_ROBId; // @[ReservationStation.scala 85:22]
  reg [3:0] entries_1_opr1; // @[ReservationStation.scala 85:22]
  reg [3:0] entries_1_opr2; // @[ReservationStation.scala 85:22]
  reg [4:0] entries_1_rs1; // @[ReservationStation.scala 85:22]
  reg [4:0] entries_1_rs2; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_1_rs1Val; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_1_rs2Val; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_1_rs1ROBId; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_1_rs2ROBId; // @[ReservationStation.scala 85:22]
  reg [2:0] entries_1_immSrc; // @[ReservationStation.scala 85:22]
  reg  entries_1_immSign; // @[ReservationStation.scala 85:22]
  reg [3:0] entries_1_excpType; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_1_pc; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_1_inst; // @[ReservationStation.scala 85:22]
  reg  entries_2_busy; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_2_op; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_2_ROBId; // @[ReservationStation.scala 85:22]
  reg [3:0] entries_2_opr1; // @[ReservationStation.scala 85:22]
  reg [3:0] entries_2_opr2; // @[ReservationStation.scala 85:22]
  reg [4:0] entries_2_rs1; // @[ReservationStation.scala 85:22]
  reg [4:0] entries_2_rs2; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_2_rs1Val; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_2_rs2Val; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_2_rs1ROBId; // @[ReservationStation.scala 85:22]
  reg [7:0] entries_2_rs2ROBId; // @[ReservationStation.scala 85:22]
  reg [2:0] entries_2_immSrc; // @[ReservationStation.scala 85:22]
  reg  entries_2_immSign; // @[ReservationStation.scala 85:22]
  reg [3:0] entries_2_excpType; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_2_pc; // @[ReservationStation.scala 85:22]
  reg [31:0] entries_2_inst; // @[ReservationStation.scala 85:22]
  reg [1:0] head; // @[ReservationStation.scala 86:23]
  reg [1:0] tail; // @[ReservationStation.scala 87:23]
  reg [1:0] count; // @[ReservationStation.scala 89:24]
  wire  full = count == 2'h3; // @[ReservationStation.scala 90:22]
  wire [7:0] _GEN_1 = 2'h1 == head ? entries_1_rs1ROBId : entries_0_rs1ROBId; // @[ReservationStation.scala 94:{41,41}]
  wire [7:0] _GEN_2 = 2'h2 == head ? entries_2_rs1ROBId : _GEN_1; // @[ReservationStation.scala 94:{41,41}]
  wire [7:0] _GEN_4 = 2'h1 == head ? entries_1_rs2ROBId : entries_0_rs2ROBId; // @[ReservationStation.scala 94:{73,73}]
  wire [7:0] _GEN_5 = 2'h2 == head ? entries_2_rs2ROBId : _GEN_4; // @[ReservationStation.scala 94:{73,73}]
  wire  oprReady = _GEN_2 == 8'h0 & _GEN_5 == 8'h0; // @[ReservationStation.scala 94:49]
  wire  _GEN_7 = 2'h1 == tail ? entries_1_busy : entries_0_busy; // @[ReservationStation.scala 95:{30,30}]
  wire  _GEN_8 = 2'h2 == tail ? entries_2_busy : _GEN_7; // @[ReservationStation.scala 95:{30,30}]
  wire  _GEN_10 = 2'h1 == head ? entries_1_busy : entries_0_busy; // @[ReservationStation.scala 96:{30,30}]
  wire  _GEN_11 = 2'h2 == head ? entries_2_busy : _GEN_10; // @[ReservationStation.scala 96:{30,30}]
  wire [7:0] _GEN_13 = 2'h1 == head ? entries_1_op : entries_0_op; // @[ReservationStation.scala 97:{20,20}]
  wire [7:0] _GEN_16 = 2'h1 == head ? entries_1_ROBId : entries_0_ROBId; // @[ReservationStation.scala 98:{23,23}]
  wire [7:0] _GEN_17 = 2'h2 == head ? entries_2_ROBId : _GEN_16; // @[ReservationStation.scala 98:{23,23}]
  wire [3:0] _GEN_19 = 2'h1 == head ? entries_1_opr1 : entries_0_opr1; // @[ReservationStation.scala 99:{22,22}]
  wire [3:0] _GEN_22 = 2'h1 == head ? entries_1_opr2 : entries_0_opr2; // @[ReservationStation.scala 100:{22,22}]
  wire [31:0] _GEN_25 = 2'h1 == head ? entries_1_rs1Val : entries_0_rs1Val; // @[ReservationStation.scala 101:{24,24}]
  wire [31:0] _GEN_28 = 2'h1 == head ? entries_1_rs2Val : entries_0_rs2Val; // @[ReservationStation.scala 102:{24,24}]
  wire [2:0] _GEN_31 = 2'h1 == head ? entries_1_immSrc : entries_0_immSrc; // @[ReservationStation.scala 103:{24,24}]
  wire  _GEN_34 = 2'h1 == head ? entries_1_immSign : entries_0_immSign; // @[ReservationStation.scala 104:{25,25}]
  wire [3:0] _GEN_37 = 2'h1 == head ? entries_1_excpType : entries_0_excpType; // @[ReservationStation.scala 105:{26,26}]
  wire [31:0] _GEN_40 = 2'h1 == head ? entries_1_pc : entries_0_pc; // @[ReservationStation.scala 106:{20,20}]
  wire [31:0] _GEN_43 = 2'h1 == head ? entries_1_inst : entries_0_inst; // @[ReservationStation.scala 107:{22,22}]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_45 = 2'h0 == tail | entries_0_busy; // @[ReservationStation.scala 121:{28,28} 85:22]
  wire  _GEN_46 = 2'h1 == tail | entries_1_busy; // @[ReservationStation.scala 121:{28,28} 85:22]
  wire  _GEN_47 = 2'h2 == tail | entries_2_busy; // @[ReservationStation.scala 121:{28,28} 85:22]
  wire [7:0] _GEN_54 = 2'h0 == tail ? io_enq_bits_rs1ROBId : entries_0_rs1ROBId; // @[ReservationStation.scala 124:{32,32} 85:22]
  wire [7:0] _GEN_55 = 2'h1 == tail ? io_enq_bits_rs1ROBId : entries_1_rs1ROBId; // @[ReservationStation.scala 124:{32,32} 85:22]
  wire [7:0] _GEN_56 = 2'h2 == tail ? io_enq_bits_rs1ROBId : entries_2_rs1ROBId; // @[ReservationStation.scala 124:{32,32} 85:22]
  wire [7:0] _GEN_57 = 2'h0 == tail ? io_enq_bits_rs2ROBId : entries_0_rs2ROBId; // @[ReservationStation.scala 125:{32,32} 85:22]
  wire [7:0] _GEN_58 = 2'h1 == tail ? io_enq_bits_rs2ROBId : entries_1_rs2ROBId; // @[ReservationStation.scala 125:{32,32} 85:22]
  wire [7:0] _GEN_59 = 2'h2 == tail ? io_enq_bits_rs2ROBId : entries_2_rs2ROBId; // @[ReservationStation.scala 125:{32,32} 85:22]
  wire [7:0] _GEN_97 = 5'h1 == io_enq_bits_rs1 ? io_regStatus_1_owner : io_regStatus_0_owner; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_98 = 5'h2 == io_enq_bits_rs1 ? io_regStatus_2_owner : _GEN_97; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_99 = 5'h3 == io_enq_bits_rs1 ? io_regStatus_3_owner : _GEN_98; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_100 = 5'h4 == io_enq_bits_rs1 ? io_regStatus_4_owner : _GEN_99; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_101 = 5'h5 == io_enq_bits_rs1 ? io_regStatus_5_owner : _GEN_100; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_102 = 5'h6 == io_enq_bits_rs1 ? io_regStatus_6_owner : _GEN_101; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_103 = 5'h7 == io_enq_bits_rs1 ? io_regStatus_7_owner : _GEN_102; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_104 = 5'h8 == io_enq_bits_rs1 ? io_regStatus_8_owner : _GEN_103; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_105 = 5'h9 == io_enq_bits_rs1 ? io_regStatus_9_owner : _GEN_104; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_106 = 5'ha == io_enq_bits_rs1 ? io_regStatus_10_owner : _GEN_105; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_107 = 5'hb == io_enq_bits_rs1 ? io_regStatus_11_owner : _GEN_106; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_108 = 5'hc == io_enq_bits_rs1 ? io_regStatus_12_owner : _GEN_107; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_109 = 5'hd == io_enq_bits_rs1 ? io_regStatus_13_owner : _GEN_108; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_110 = 5'he == io_enq_bits_rs1 ? io_regStatus_14_owner : _GEN_109; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_111 = 5'hf == io_enq_bits_rs1 ? io_regStatus_15_owner : _GEN_110; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_112 = 5'h10 == io_enq_bits_rs1 ? io_regStatus_16_owner : _GEN_111; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_113 = 5'h11 == io_enq_bits_rs1 ? io_regStatus_17_owner : _GEN_112; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_114 = 5'h12 == io_enq_bits_rs1 ? io_regStatus_18_owner : _GEN_113; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_115 = 5'h13 == io_enq_bits_rs1 ? io_regStatus_19_owner : _GEN_114; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_116 = 5'h14 == io_enq_bits_rs1 ? io_regStatus_20_owner : _GEN_115; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_117 = 5'h15 == io_enq_bits_rs1 ? io_regStatus_21_owner : _GEN_116; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_118 = 5'h16 == io_enq_bits_rs1 ? io_regStatus_22_owner : _GEN_117; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_119 = 5'h17 == io_enq_bits_rs1 ? io_regStatus_23_owner : _GEN_118; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_120 = 5'h18 == io_enq_bits_rs1 ? io_regStatus_24_owner : _GEN_119; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_121 = 5'h19 == io_enq_bits_rs1 ? io_regStatus_25_owner : _GEN_120; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_122 = 5'h1a == io_enq_bits_rs1 ? io_regStatus_26_owner : _GEN_121; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_123 = 5'h1b == io_enq_bits_rs1 ? io_regStatus_27_owner : _GEN_122; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_124 = 5'h1c == io_enq_bits_rs1 ? io_regStatus_28_owner : _GEN_123; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_125 = 5'h1d == io_enq_bits_rs1 ? io_regStatus_29_owner : _GEN_124; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_126 = 5'h1e == io_enq_bits_rs1 ? io_regStatus_30_owner : _GEN_125; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_127 = 5'h1f == io_enq_bits_rs1 ? io_regStatus_31_owner : _GEN_126; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_93 = 2'h0 == tail ? _GEN_127 : _GEN_54; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_94 = 2'h1 == tail ? _GEN_127 : _GEN_55; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_95 = 2'h2 == tail ? _GEN_127 : _GEN_56; // @[ReservationStation.scala 140:{32,32}]
  wire [7:0] _GEN_132 = 5'h1 == io_enq_bits_rs2 ? io_regStatus_1_owner : io_regStatus_0_owner; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_133 = 5'h2 == io_enq_bits_rs2 ? io_regStatus_2_owner : _GEN_132; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_134 = 5'h3 == io_enq_bits_rs2 ? io_regStatus_3_owner : _GEN_133; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_135 = 5'h4 == io_enq_bits_rs2 ? io_regStatus_4_owner : _GEN_134; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_136 = 5'h5 == io_enq_bits_rs2 ? io_regStatus_5_owner : _GEN_135; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_137 = 5'h6 == io_enq_bits_rs2 ? io_regStatus_6_owner : _GEN_136; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_138 = 5'h7 == io_enq_bits_rs2 ? io_regStatus_7_owner : _GEN_137; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_139 = 5'h8 == io_enq_bits_rs2 ? io_regStatus_8_owner : _GEN_138; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_140 = 5'h9 == io_enq_bits_rs2 ? io_regStatus_9_owner : _GEN_139; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_141 = 5'ha == io_enq_bits_rs2 ? io_regStatus_10_owner : _GEN_140; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_142 = 5'hb == io_enq_bits_rs2 ? io_regStatus_11_owner : _GEN_141; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_143 = 5'hc == io_enq_bits_rs2 ? io_regStatus_12_owner : _GEN_142; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_144 = 5'hd == io_enq_bits_rs2 ? io_regStatus_13_owner : _GEN_143; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_145 = 5'he == io_enq_bits_rs2 ? io_regStatus_14_owner : _GEN_144; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_146 = 5'hf == io_enq_bits_rs2 ? io_regStatus_15_owner : _GEN_145; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_147 = 5'h10 == io_enq_bits_rs2 ? io_regStatus_16_owner : _GEN_146; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_148 = 5'h11 == io_enq_bits_rs2 ? io_regStatus_17_owner : _GEN_147; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_149 = 5'h12 == io_enq_bits_rs2 ? io_regStatus_18_owner : _GEN_148; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_150 = 5'h13 == io_enq_bits_rs2 ? io_regStatus_19_owner : _GEN_149; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_151 = 5'h14 == io_enq_bits_rs2 ? io_regStatus_20_owner : _GEN_150; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_152 = 5'h15 == io_enq_bits_rs2 ? io_regStatus_21_owner : _GEN_151; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_153 = 5'h16 == io_enq_bits_rs2 ? io_regStatus_22_owner : _GEN_152; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_154 = 5'h17 == io_enq_bits_rs2 ? io_regStatus_23_owner : _GEN_153; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_155 = 5'h18 == io_enq_bits_rs2 ? io_regStatus_24_owner : _GEN_154; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_156 = 5'h19 == io_enq_bits_rs2 ? io_regStatus_25_owner : _GEN_155; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_157 = 5'h1a == io_enq_bits_rs2 ? io_regStatus_26_owner : _GEN_156; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_158 = 5'h1b == io_enq_bits_rs2 ? io_regStatus_27_owner : _GEN_157; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_159 = 5'h1c == io_enq_bits_rs2 ? io_regStatus_28_owner : _GEN_158; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_160 = 5'h1d == io_enq_bits_rs2 ? io_regStatus_29_owner : _GEN_159; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_161 = 5'h1e == io_enq_bits_rs2 ? io_regStatus_30_owner : _GEN_160; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_162 = 5'h1f == io_enq_bits_rs2 ? io_regStatus_31_owner : _GEN_161; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_128 = 2'h0 == tail ? _GEN_162 : _GEN_57; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_129 = 2'h1 == tail ? _GEN_162 : _GEN_58; // @[ReservationStation.scala 141:{32,32}]
  wire [7:0] _GEN_130 = 2'h2 == tail ? _GEN_162 : _GEN_59; // @[ReservationStation.scala 141:{32,32}]
  wire [31:0] _GEN_163 = 2'h0 == tail ? io_rf_0_data : entries_0_rs1Val; // @[ReservationStation.scala 146:{30,30} 85:22]
  wire [31:0] _GEN_164 = 2'h1 == tail ? io_rf_0_data : entries_1_rs1Val; // @[ReservationStation.scala 146:{30,30} 85:22]
  wire [31:0] _GEN_165 = 2'h2 == tail ? io_rf_0_data : entries_2_rs1Val; // @[ReservationStation.scala 146:{30,30} 85:22]
  wire [31:0] _GEN_166 = 2'h0 == tail ? io_rf_1_data : entries_0_rs2Val; // @[ReservationStation.scala 147:{30,30} 85:22]
  wire [31:0] _GEN_167 = 2'h1 == tail ? io_rf_1_data : entries_1_rs2Val; // @[ReservationStation.scala 147:{30,30} 85:22]
  wire [31:0] _GEN_168 = 2'h2 == tail ? io_rf_1_data : entries_2_rs2Val; // @[ReservationStation.scala 147:{30,30} 85:22]
  wire [1:0] _tail_T_2 = tail + 2'h1; // @[ReservationStation.scala 149:60]
  wire  _GEN_169 = _T ? _GEN_45 : entries_0_busy; // @[ReservationStation.scala 120:24 85:22]
  wire  _GEN_170 = _T ? _GEN_46 : entries_1_busy; // @[ReservationStation.scala 120:24 85:22]
  wire  _GEN_171 = _T ? _GEN_47 : entries_2_busy; // @[ReservationStation.scala 120:24 85:22]
  wire [7:0] _GEN_178 = _T ? _GEN_93 : entries_0_rs1ROBId; // @[ReservationStation.scala 120:24 85:22]
  wire [7:0] _GEN_179 = _T ? _GEN_94 : entries_1_rs1ROBId; // @[ReservationStation.scala 120:24 85:22]
  wire [7:0] _GEN_180 = _T ? _GEN_95 : entries_2_rs1ROBId; // @[ReservationStation.scala 120:24 85:22]
  wire [7:0] _GEN_181 = _T ? _GEN_128 : entries_0_rs2ROBId; // @[ReservationStation.scala 120:24 85:22]
  wire [7:0] _GEN_182 = _T ? _GEN_129 : entries_1_rs2ROBId; // @[ReservationStation.scala 120:24 85:22]
  wire [7:0] _GEN_183 = _T ? _GEN_130 : entries_2_rs2ROBId; // @[ReservationStation.scala 120:24 85:22]
  wire [31:0] _GEN_216 = _T ? _GEN_163 : entries_0_rs1Val; // @[ReservationStation.scala 120:24 85:22]
  wire [31:0] _GEN_217 = _T ? _GEN_164 : entries_1_rs1Val; // @[ReservationStation.scala 120:24 85:22]
  wire [31:0] _GEN_218 = _T ? _GEN_165 : entries_2_rs1Val; // @[ReservationStation.scala 120:24 85:22]
  wire [31:0] _GEN_219 = _T ? _GEN_166 : entries_0_rs2Val; // @[ReservationStation.scala 120:24 85:22]
  wire [31:0] _GEN_220 = _T ? _GEN_167 : entries_1_rs2Val; // @[ReservationStation.scala 120:24 85:22]
  wire [31:0] _GEN_221 = _T ? _GEN_168 : entries_2_rs2Val; // @[ReservationStation.scala 120:24 85:22]
  wire  _T_1 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _head_T_2 = head + 2'h1; // @[ReservationStation.scala 158:60]
  wire [7:0] _GEN_233 = _T_1 ? _GEN_17 : 8'h0; // @[ReservationStation.scala 110:23 152:24 155:27]
  wire [1:0] _count_T_1 = count + 2'h1; // @[ReservationStation.scala 163:28]
  wire [1:0] _GEN_236 = _T ? _count_T_1 : count; // @[ReservationStation.scala 162:27 163:19 89:24]
  wire [1:0] _count_T_3 = count - 2'h1; // @[ReservationStation.scala 166:28]
  wire [7:0] _rs1ROBEntry_T_1 = entries_0_rs1ROBId - 8'h1; // @[ReservationStation.scala 178:53]
  wire [7:0] _rs2ROBEntry_T_1 = entries_0_rs2ROBId - 8'h1; // @[ReservationStation.scala 179:53]
  wire [1:0] _GEN_240 = 3'h1 == _rs1ROBEntry_T_1[2:0] ? io_robRead_1_state : io_robRead_0_state; // @[ReservationStation.scala 180:{69,69}]
  wire [1:0] _GEN_241 = 3'h2 == _rs1ROBEntry_T_1[2:0] ? io_robRead_2_state : _GEN_240; // @[ReservationStation.scala 180:{69,69}]
  wire [1:0] _GEN_242 = 3'h3 == _rs1ROBEntry_T_1[2:0] ? io_robRead_3_state : _GEN_241; // @[ReservationStation.scala 180:{69,69}]
  wire [1:0] _GEN_243 = 3'h4 == _rs1ROBEntry_T_1[2:0] ? io_robRead_4_state : _GEN_242; // @[ReservationStation.scala 180:{69,69}]
  wire  _GEN_245 = 3'h1 == _rs1ROBEntry_T_1[2:0] ? io_robRead_1_busy : io_robRead_0_busy; // @[ReservationStation.scala 180:{48,48}]
  wire  _GEN_246 = 3'h2 == _rs1ROBEntry_T_1[2:0] ? io_robRead_2_busy : _GEN_245; // @[ReservationStation.scala 180:{48,48}]
  wire  _GEN_247 = 3'h3 == _rs1ROBEntry_T_1[2:0] ? io_robRead_3_busy : _GEN_246; // @[ReservationStation.scala 180:{48,48}]
  wire  _GEN_248 = 3'h4 == _rs1ROBEntry_T_1[2:0] ? io_robRead_4_busy : _GEN_247; // @[ReservationStation.scala 180:{48,48}]
  wire [4:0] _GEN_250 = 3'h1 == _rs1ROBEntry_T_1[2:0] ? io_robRead_1_rd : io_robRead_0_rd; // @[ReservationStation.scala 180:{132,132}]
  wire [4:0] _GEN_251 = 3'h2 == _rs1ROBEntry_T_1[2:0] ? io_robRead_2_rd : _GEN_250; // @[ReservationStation.scala 180:{132,132}]
  wire [4:0] _GEN_252 = 3'h3 == _rs1ROBEntry_T_1[2:0] ? io_robRead_3_rd : _GEN_251; // @[ReservationStation.scala 180:{132,132}]
  wire [4:0] _GEN_253 = 3'h4 == _rs1ROBEntry_T_1[2:0] ? io_robRead_4_rd : _GEN_252; // @[ReservationStation.scala 180:{132,132}]
  wire  rs1FromROB = (_GEN_248 & _GEN_243 == 2'h2 | _GEN_243 == 2'h3) & _GEN_253 == entries_0_rs1 & entries_0_rs1 != 5'h0
    ; // @[ReservationStation.scala 180:142]
  wire [1:0] _GEN_255 = 3'h1 == _rs2ROBEntry_T_1[2:0] ? io_robRead_1_state : io_robRead_0_state; // @[ReservationStation.scala 181:{69,69}]
  wire [1:0] _GEN_256 = 3'h2 == _rs2ROBEntry_T_1[2:0] ? io_robRead_2_state : _GEN_255; // @[ReservationStation.scala 181:{69,69}]
  wire [1:0] _GEN_257 = 3'h3 == _rs2ROBEntry_T_1[2:0] ? io_robRead_3_state : _GEN_256; // @[ReservationStation.scala 181:{69,69}]
  wire [1:0] _GEN_258 = 3'h4 == _rs2ROBEntry_T_1[2:0] ? io_robRead_4_state : _GEN_257; // @[ReservationStation.scala 181:{69,69}]
  wire  _GEN_260 = 3'h1 == _rs2ROBEntry_T_1[2:0] ? io_robRead_1_busy : io_robRead_0_busy; // @[ReservationStation.scala 181:{48,48}]
  wire  _GEN_261 = 3'h2 == _rs2ROBEntry_T_1[2:0] ? io_robRead_2_busy : _GEN_260; // @[ReservationStation.scala 181:{48,48}]
  wire  _GEN_262 = 3'h3 == _rs2ROBEntry_T_1[2:0] ? io_robRead_3_busy : _GEN_261; // @[ReservationStation.scala 181:{48,48}]
  wire  _GEN_263 = 3'h4 == _rs2ROBEntry_T_1[2:0] ? io_robRead_4_busy : _GEN_262; // @[ReservationStation.scala 181:{48,48}]
  wire [4:0] _GEN_265 = 3'h1 == _rs2ROBEntry_T_1[2:0] ? io_robRead_1_rd : io_robRead_0_rd; // @[ReservationStation.scala 181:{132,132}]
  wire [4:0] _GEN_266 = 3'h2 == _rs2ROBEntry_T_1[2:0] ? io_robRead_2_rd : _GEN_265; // @[ReservationStation.scala 181:{132,132}]
  wire [4:0] _GEN_267 = 3'h3 == _rs2ROBEntry_T_1[2:0] ? io_robRead_3_rd : _GEN_266; // @[ReservationStation.scala 181:{132,132}]
  wire [4:0] _GEN_268 = 3'h4 == _rs2ROBEntry_T_1[2:0] ? io_robRead_4_rd : _GEN_267; // @[ReservationStation.scala 181:{132,132}]
  wire  rs2FromROB = (_GEN_263 & _GEN_258 == 2'h2 | _GEN_258 == 2'h3) & _GEN_268 == entries_0_rs2 & entries_0_rs2 != 5'h0
    ; // @[ReservationStation.scala 181:142]
  wire  _T_8 = entries_0_rs1ROBId != 8'h0; // @[ReservationStation.scala 182:43]
  wire [31:0] _GEN_270 = 3'h1 == _rs1ROBEntry_T_1[2:0] ? io_robRead_1_data : io_robRead_0_data; // @[ReservationStation.scala 183:{26,26}]
  wire [31:0] _GEN_271 = 3'h2 == _rs1ROBEntry_T_1[2:0] ? io_robRead_2_data : _GEN_270; // @[ReservationStation.scala 183:{26,26}]
  wire [31:0] _GEN_272 = 3'h3 == _rs1ROBEntry_T_1[2:0] ? io_robRead_3_data : _GEN_271; // @[ReservationStation.scala 183:{26,26}]
  wire  _T_10 = entries_0_rs2ROBId != 8'h0; // @[ReservationStation.scala 186:43]
  wire [31:0] _GEN_277 = 3'h1 == _rs2ROBEntry_T_1[2:0] ? io_robRead_1_data : io_robRead_0_data; // @[ReservationStation.scala 187:{26,26}]
  wire [31:0] _GEN_278 = 3'h2 == _rs2ROBEntry_T_1[2:0] ? io_robRead_2_data : _GEN_277; // @[ReservationStation.scala 187:{26,26}]
  wire [31:0] _GEN_279 = 3'h3 == _rs2ROBEntry_T_1[2:0] ? io_robRead_3_data : _GEN_278; // @[ReservationStation.scala 187:{26,26}]
  wire  _rs1MatchVec_T = io_cdb_0_bits_rd == entries_0_rs1; // @[ReservationStation.scala 192:61]
  wire  _rs1MatchVec_T_1 = io_cdb_1_bits_rd == entries_0_rs1; // @[ReservationStation.scala 192:61]
  wire  _rs1MatchVec_T_2 = io_cdb_2_bits_rd == entries_0_rs1; // @[ReservationStation.scala 192:61]
  wire  _rs1MatchVec_T_3 = io_cdb_3_bits_rd == entries_0_rs1; // @[ReservationStation.scala 192:61]
  wire [3:0] rs1MatchVec = {_rs1MatchVec_T_3,_rs1MatchVec_T_2,_rs1MatchVec_T_1,_rs1MatchVec_T}; // @[Cat.scala 33:92]
  wire  _rs2MatchVec_T = io_cdb_0_bits_rd == entries_0_rs2; // @[ReservationStation.scala 193:61]
  wire  _rs2MatchVec_T_1 = io_cdb_1_bits_rd == entries_0_rs2; // @[ReservationStation.scala 193:61]
  wire  _rs2MatchVec_T_2 = io_cdb_2_bits_rd == entries_0_rs2; // @[ReservationStation.scala 193:61]
  wire  _rs2MatchVec_T_3 = io_cdb_3_bits_rd == entries_0_rs2; // @[ReservationStation.scala 193:61]
  wire [3:0] rs2MatchVec = {_rs2MatchVec_T_3,_rs2MatchVec_T_2,_rs2MatchVec_T_1,_rs2MatchVec_T}; // @[Cat.scala 33:92]
  wire  _rs1IDMatchVec_T = io_cdb_0_bits_id == entries_0_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire  _rs1IDMatchVec_T_1 = io_cdb_1_bits_id == entries_0_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire  _rs1IDMatchVec_T_2 = io_cdb_2_bits_id == entries_0_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire  _rs1IDMatchVec_T_3 = io_cdb_3_bits_id == entries_0_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire [3:0] rs1IDMatchVec = {_rs1IDMatchVec_T_3,_rs1IDMatchVec_T_2,_rs1IDMatchVec_T_1,_rs1IDMatchVec_T}; // @[Cat.scala 33:92]
  wire  _rs2IDMatchVec_T = io_cdb_0_bits_id == entries_0_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire  _rs2IDMatchVec_T_1 = io_cdb_1_bits_id == entries_0_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire  _rs2IDMatchVec_T_2 = io_cdb_2_bits_id == entries_0_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire  _rs2IDMatchVec_T_3 = io_cdb_3_bits_id == entries_0_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire [3:0] rs2IDMatchVec = {_rs2IDMatchVec_T_3,_rs2IDMatchVec_T_2,_rs2IDMatchVec_T_1,_rs2IDMatchVec_T}; // @[Cat.scala 33:92]
  wire [3:0] cdbValidVec = {io_cdb_3_valid,io_cdb_2_valid,io_cdb_1_valid,io_cdb_0_valid}; // @[Cat.scala 33:92]
  wire [3:0] _cdbBypassRs1_T = cdbValidVec & rs1MatchVec; // @[ReservationStation.scala 197:44]
  wire [3:0] cdbBypassRs1 = _cdbBypassRs1_T & rs1IDMatchVec; // @[ReservationStation.scala 197:58]
  wire [3:0] _cdbBypassRs2_T = cdbValidVec & rs2MatchVec; // @[ReservationStation.scala 198:44]
  wire [3:0] cdbBypassRs2 = _cdbBypassRs2_T & rs2IDMatchVec; // @[ReservationStation.scala 198:58]
  wire  bypassRs1 = |cdbBypassRs1; // @[ReservationStation.scala 200:42]
  wire  bypassRs2 = |cdbBypassRs2; // @[ReservationStation.scala 201:42]
  wire [31:0] _entries_0_rs1Val_T_4 = cdbBypassRs1[0] ? io_cdb_0_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs1Val_T_5 = cdbBypassRs1[1] ? io_cdb_1_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs1Val_T_6 = cdbBypassRs1[2] ? io_cdb_2_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs1Val_T_7 = cdbBypassRs1[3] ? io_cdb_3_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs1Val_T_8 = _entries_0_rs1Val_T_4 | _entries_0_rs1Val_T_5; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs1Val_T_9 = _entries_0_rs1Val_T_8 | _entries_0_rs1Val_T_6; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs1Val_T_10 = _entries_0_rs1Val_T_9 | _entries_0_rs1Val_T_7; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs2Val_T_4 = cdbBypassRs2[0] ? io_cdb_0_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs2Val_T_5 = cdbBypassRs2[1] ? io_cdb_1_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs2Val_T_6 = cdbBypassRs2[2] ? io_cdb_2_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs2Val_T_7 = cdbBypassRs2[3] ? io_cdb_3_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs2Val_T_8 = _entries_0_rs2Val_T_4 | _entries_0_rs2Val_T_5; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs2Val_T_9 = _entries_0_rs2Val_T_8 | _entries_0_rs2Val_T_6; // @[Mux.scala 27:73]
  wire [31:0] _entries_0_rs2Val_T_10 = _entries_0_rs2Val_T_9 | _entries_0_rs2Val_T_7; // @[Mux.scala 27:73]
  wire [7:0] _rs1ROBEntry_T_4 = entries_1_rs1ROBId - 8'h1; // @[ReservationStation.scala 178:53]
  wire [7:0] _rs2ROBEntry_T_4 = entries_1_rs2ROBId - 8'h1; // @[ReservationStation.scala 179:53]
  wire [1:0] _GEN_292 = 3'h1 == _rs1ROBEntry_T_4[2:0] ? io_robRead_1_state : io_robRead_0_state; // @[ReservationStation.scala 180:{69,69}]
  wire [1:0] _GEN_293 = 3'h2 == _rs1ROBEntry_T_4[2:0] ? io_robRead_2_state : _GEN_292; // @[ReservationStation.scala 180:{69,69}]
  wire [1:0] _GEN_294 = 3'h3 == _rs1ROBEntry_T_4[2:0] ? io_robRead_3_state : _GEN_293; // @[ReservationStation.scala 180:{69,69}]
  wire [1:0] _GEN_295 = 3'h4 == _rs1ROBEntry_T_4[2:0] ? io_robRead_4_state : _GEN_294; // @[ReservationStation.scala 180:{69,69}]
  wire  _GEN_297 = 3'h1 == _rs1ROBEntry_T_4[2:0] ? io_robRead_1_busy : io_robRead_0_busy; // @[ReservationStation.scala 180:{48,48}]
  wire  _GEN_298 = 3'h2 == _rs1ROBEntry_T_4[2:0] ? io_robRead_2_busy : _GEN_297; // @[ReservationStation.scala 180:{48,48}]
  wire  _GEN_299 = 3'h3 == _rs1ROBEntry_T_4[2:0] ? io_robRead_3_busy : _GEN_298; // @[ReservationStation.scala 180:{48,48}]
  wire  _GEN_300 = 3'h4 == _rs1ROBEntry_T_4[2:0] ? io_robRead_4_busy : _GEN_299; // @[ReservationStation.scala 180:{48,48}]
  wire [4:0] _GEN_302 = 3'h1 == _rs1ROBEntry_T_4[2:0] ? io_robRead_1_rd : io_robRead_0_rd; // @[ReservationStation.scala 180:{132,132}]
  wire [4:0] _GEN_303 = 3'h2 == _rs1ROBEntry_T_4[2:0] ? io_robRead_2_rd : _GEN_302; // @[ReservationStation.scala 180:{132,132}]
  wire [4:0] _GEN_304 = 3'h3 == _rs1ROBEntry_T_4[2:0] ? io_robRead_3_rd : _GEN_303; // @[ReservationStation.scala 180:{132,132}]
  wire [4:0] _GEN_305 = 3'h4 == _rs1ROBEntry_T_4[2:0] ? io_robRead_4_rd : _GEN_304; // @[ReservationStation.scala 180:{132,132}]
  wire  rs1FromROB_1 = (_GEN_300 & _GEN_295 == 2'h2 | _GEN_295 == 2'h3) & _GEN_305 == entries_1_rs1 & entries_1_rs1 != 5'h0
    ; // @[ReservationStation.scala 180:142]
  wire [1:0] _GEN_307 = 3'h1 == _rs2ROBEntry_T_4[2:0] ? io_robRead_1_state : io_robRead_0_state; // @[ReservationStation.scala 181:{69,69}]
  wire [1:0] _GEN_308 = 3'h2 == _rs2ROBEntry_T_4[2:0] ? io_robRead_2_state : _GEN_307; // @[ReservationStation.scala 181:{69,69}]
  wire [1:0] _GEN_309 = 3'h3 == _rs2ROBEntry_T_4[2:0] ? io_robRead_3_state : _GEN_308; // @[ReservationStation.scala 181:{69,69}]
  wire [1:0] _GEN_310 = 3'h4 == _rs2ROBEntry_T_4[2:0] ? io_robRead_4_state : _GEN_309; // @[ReservationStation.scala 181:{69,69}]
  wire  _GEN_312 = 3'h1 == _rs2ROBEntry_T_4[2:0] ? io_robRead_1_busy : io_robRead_0_busy; // @[ReservationStation.scala 181:{48,48}]
  wire  _GEN_313 = 3'h2 == _rs2ROBEntry_T_4[2:0] ? io_robRead_2_busy : _GEN_312; // @[ReservationStation.scala 181:{48,48}]
  wire  _GEN_314 = 3'h3 == _rs2ROBEntry_T_4[2:0] ? io_robRead_3_busy : _GEN_313; // @[ReservationStation.scala 181:{48,48}]
  wire  _GEN_315 = 3'h4 == _rs2ROBEntry_T_4[2:0] ? io_robRead_4_busy : _GEN_314; // @[ReservationStation.scala 181:{48,48}]
  wire [4:0] _GEN_317 = 3'h1 == _rs2ROBEntry_T_4[2:0] ? io_robRead_1_rd : io_robRead_0_rd; // @[ReservationStation.scala 181:{132,132}]
  wire [4:0] _GEN_318 = 3'h2 == _rs2ROBEntry_T_4[2:0] ? io_robRead_2_rd : _GEN_317; // @[ReservationStation.scala 181:{132,132}]
  wire [4:0] _GEN_319 = 3'h3 == _rs2ROBEntry_T_4[2:0] ? io_robRead_3_rd : _GEN_318; // @[ReservationStation.scala 181:{132,132}]
  wire [4:0] _GEN_320 = 3'h4 == _rs2ROBEntry_T_4[2:0] ? io_robRead_4_rd : _GEN_319; // @[ReservationStation.scala 181:{132,132}]
  wire  rs2FromROB_1 = (_GEN_315 & _GEN_310 == 2'h2 | _GEN_310 == 2'h3) & _GEN_320 == entries_1_rs2 & entries_1_rs2 != 5'h0
    ; // @[ReservationStation.scala 181:142]
  wire  _T_16 = entries_1_rs1ROBId != 8'h0; // @[ReservationStation.scala 182:43]
  wire [31:0] _GEN_322 = 3'h1 == _rs1ROBEntry_T_4[2:0] ? io_robRead_1_data : io_robRead_0_data; // @[ReservationStation.scala 183:{26,26}]
  wire [31:0] _GEN_323 = 3'h2 == _rs1ROBEntry_T_4[2:0] ? io_robRead_2_data : _GEN_322; // @[ReservationStation.scala 183:{26,26}]
  wire [31:0] _GEN_324 = 3'h3 == _rs1ROBEntry_T_4[2:0] ? io_robRead_3_data : _GEN_323; // @[ReservationStation.scala 183:{26,26}]
  wire  _T_18 = entries_1_rs2ROBId != 8'h0; // @[ReservationStation.scala 186:43]
  wire [31:0] _GEN_329 = 3'h1 == _rs2ROBEntry_T_4[2:0] ? io_robRead_1_data : io_robRead_0_data; // @[ReservationStation.scala 187:{26,26}]
  wire [31:0] _GEN_330 = 3'h2 == _rs2ROBEntry_T_4[2:0] ? io_robRead_2_data : _GEN_329; // @[ReservationStation.scala 187:{26,26}]
  wire [31:0] _GEN_331 = 3'h3 == _rs2ROBEntry_T_4[2:0] ? io_robRead_3_data : _GEN_330; // @[ReservationStation.scala 187:{26,26}]
  wire  _rs1MatchVec_T_4 = io_cdb_0_bits_rd == entries_1_rs1; // @[ReservationStation.scala 192:61]
  wire  _rs1MatchVec_T_5 = io_cdb_1_bits_rd == entries_1_rs1; // @[ReservationStation.scala 192:61]
  wire  _rs1MatchVec_T_6 = io_cdb_2_bits_rd == entries_1_rs1; // @[ReservationStation.scala 192:61]
  wire  _rs1MatchVec_T_7 = io_cdb_3_bits_rd == entries_1_rs1; // @[ReservationStation.scala 192:61]
  wire [3:0] rs1MatchVec_1 = {_rs1MatchVec_T_7,_rs1MatchVec_T_6,_rs1MatchVec_T_5,_rs1MatchVec_T_4}; // @[Cat.scala 33:92]
  wire  _rs2MatchVec_T_4 = io_cdb_0_bits_rd == entries_1_rs2; // @[ReservationStation.scala 193:61]
  wire  _rs2MatchVec_T_5 = io_cdb_1_bits_rd == entries_1_rs2; // @[ReservationStation.scala 193:61]
  wire  _rs2MatchVec_T_6 = io_cdb_2_bits_rd == entries_1_rs2; // @[ReservationStation.scala 193:61]
  wire  _rs2MatchVec_T_7 = io_cdb_3_bits_rd == entries_1_rs2; // @[ReservationStation.scala 193:61]
  wire [3:0] rs2MatchVec_1 = {_rs2MatchVec_T_7,_rs2MatchVec_T_6,_rs2MatchVec_T_5,_rs2MatchVec_T_4}; // @[Cat.scala 33:92]
  wire  _rs1IDMatchVec_T_4 = io_cdb_0_bits_id == entries_1_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire  _rs1IDMatchVec_T_5 = io_cdb_1_bits_id == entries_1_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire  _rs1IDMatchVec_T_6 = io_cdb_2_bits_id == entries_1_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire  _rs1IDMatchVec_T_7 = io_cdb_3_bits_id == entries_1_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire [3:0] rs1IDMatchVec_1 = {_rs1IDMatchVec_T_7,_rs1IDMatchVec_T_6,_rs1IDMatchVec_T_5,_rs1IDMatchVec_T_4}; // @[Cat.scala 33:92]
  wire  _rs2IDMatchVec_T_4 = io_cdb_0_bits_id == entries_1_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire  _rs2IDMatchVec_T_5 = io_cdb_1_bits_id == entries_1_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire  _rs2IDMatchVec_T_6 = io_cdb_2_bits_id == entries_1_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire  _rs2IDMatchVec_T_7 = io_cdb_3_bits_id == entries_1_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire [3:0] rs2IDMatchVec_1 = {_rs2IDMatchVec_T_7,_rs2IDMatchVec_T_6,_rs2IDMatchVec_T_5,_rs2IDMatchVec_T_4}; // @[Cat.scala 33:92]
  wire [3:0] _cdbBypassRs1_T_1 = cdbValidVec & rs1MatchVec_1; // @[ReservationStation.scala 197:44]
  wire [3:0] cdbBypassRs1_1 = _cdbBypassRs1_T_1 & rs1IDMatchVec_1; // @[ReservationStation.scala 197:58]
  wire [3:0] _cdbBypassRs2_T_1 = cdbValidVec & rs2MatchVec_1; // @[ReservationStation.scala 198:44]
  wire [3:0] cdbBypassRs2_1 = _cdbBypassRs2_T_1 & rs2IDMatchVec_1; // @[ReservationStation.scala 198:58]
  wire  bypassRs1_1 = |cdbBypassRs1_1; // @[ReservationStation.scala 200:42]
  wire  bypassRs2_1 = |cdbBypassRs2_1; // @[ReservationStation.scala 201:42]
  wire [31:0] _entries_1_rs1Val_T_4 = cdbBypassRs1_1[0] ? io_cdb_0_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs1Val_T_5 = cdbBypassRs1_1[1] ? io_cdb_1_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs1Val_T_6 = cdbBypassRs1_1[2] ? io_cdb_2_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs1Val_T_7 = cdbBypassRs1_1[3] ? io_cdb_3_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs1Val_T_8 = _entries_1_rs1Val_T_4 | _entries_1_rs1Val_T_5; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs1Val_T_9 = _entries_1_rs1Val_T_8 | _entries_1_rs1Val_T_6; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs1Val_T_10 = _entries_1_rs1Val_T_9 | _entries_1_rs1Val_T_7; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs2Val_T_4 = cdbBypassRs2_1[0] ? io_cdb_0_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs2Val_T_5 = cdbBypassRs2_1[1] ? io_cdb_1_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs2Val_T_6 = cdbBypassRs2_1[2] ? io_cdb_2_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs2Val_T_7 = cdbBypassRs2_1[3] ? io_cdb_3_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs2Val_T_8 = _entries_1_rs2Val_T_4 | _entries_1_rs2Val_T_5; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs2Val_T_9 = _entries_1_rs2Val_T_8 | _entries_1_rs2Val_T_6; // @[Mux.scala 27:73]
  wire [31:0] _entries_1_rs2Val_T_10 = _entries_1_rs2Val_T_9 | _entries_1_rs2Val_T_7; // @[Mux.scala 27:73]
  wire [7:0] _rs1ROBEntry_T_7 = entries_2_rs1ROBId - 8'h1; // @[ReservationStation.scala 178:53]
  wire [7:0] _rs2ROBEntry_T_7 = entries_2_rs2ROBId - 8'h1; // @[ReservationStation.scala 179:53]
  wire [1:0] _GEN_344 = 3'h1 == _rs1ROBEntry_T_7[2:0] ? io_robRead_1_state : io_robRead_0_state; // @[ReservationStation.scala 180:{69,69}]
  wire [1:0] _GEN_345 = 3'h2 == _rs1ROBEntry_T_7[2:0] ? io_robRead_2_state : _GEN_344; // @[ReservationStation.scala 180:{69,69}]
  wire [1:0] _GEN_346 = 3'h3 == _rs1ROBEntry_T_7[2:0] ? io_robRead_3_state : _GEN_345; // @[ReservationStation.scala 180:{69,69}]
  wire [1:0] _GEN_347 = 3'h4 == _rs1ROBEntry_T_7[2:0] ? io_robRead_4_state : _GEN_346; // @[ReservationStation.scala 180:{69,69}]
  wire  _GEN_349 = 3'h1 == _rs1ROBEntry_T_7[2:0] ? io_robRead_1_busy : io_robRead_0_busy; // @[ReservationStation.scala 180:{48,48}]
  wire  _GEN_350 = 3'h2 == _rs1ROBEntry_T_7[2:0] ? io_robRead_2_busy : _GEN_349; // @[ReservationStation.scala 180:{48,48}]
  wire  _GEN_351 = 3'h3 == _rs1ROBEntry_T_7[2:0] ? io_robRead_3_busy : _GEN_350; // @[ReservationStation.scala 180:{48,48}]
  wire  _GEN_352 = 3'h4 == _rs1ROBEntry_T_7[2:0] ? io_robRead_4_busy : _GEN_351; // @[ReservationStation.scala 180:{48,48}]
  wire [4:0] _GEN_354 = 3'h1 == _rs1ROBEntry_T_7[2:0] ? io_robRead_1_rd : io_robRead_0_rd; // @[ReservationStation.scala 180:{132,132}]
  wire [4:0] _GEN_355 = 3'h2 == _rs1ROBEntry_T_7[2:0] ? io_robRead_2_rd : _GEN_354; // @[ReservationStation.scala 180:{132,132}]
  wire [4:0] _GEN_356 = 3'h3 == _rs1ROBEntry_T_7[2:0] ? io_robRead_3_rd : _GEN_355; // @[ReservationStation.scala 180:{132,132}]
  wire [4:0] _GEN_357 = 3'h4 == _rs1ROBEntry_T_7[2:0] ? io_robRead_4_rd : _GEN_356; // @[ReservationStation.scala 180:{132,132}]
  wire  rs1FromROB_2 = (_GEN_352 & _GEN_347 == 2'h2 | _GEN_347 == 2'h3) & _GEN_357 == entries_2_rs1 & entries_2_rs1 != 5'h0
    ; // @[ReservationStation.scala 180:142]
  wire [1:0] _GEN_359 = 3'h1 == _rs2ROBEntry_T_7[2:0] ? io_robRead_1_state : io_robRead_0_state; // @[ReservationStation.scala 181:{69,69}]
  wire [1:0] _GEN_360 = 3'h2 == _rs2ROBEntry_T_7[2:0] ? io_robRead_2_state : _GEN_359; // @[ReservationStation.scala 181:{69,69}]
  wire [1:0] _GEN_361 = 3'h3 == _rs2ROBEntry_T_7[2:0] ? io_robRead_3_state : _GEN_360; // @[ReservationStation.scala 181:{69,69}]
  wire [1:0] _GEN_362 = 3'h4 == _rs2ROBEntry_T_7[2:0] ? io_robRead_4_state : _GEN_361; // @[ReservationStation.scala 181:{69,69}]
  wire  _GEN_364 = 3'h1 == _rs2ROBEntry_T_7[2:0] ? io_robRead_1_busy : io_robRead_0_busy; // @[ReservationStation.scala 181:{48,48}]
  wire  _GEN_365 = 3'h2 == _rs2ROBEntry_T_7[2:0] ? io_robRead_2_busy : _GEN_364; // @[ReservationStation.scala 181:{48,48}]
  wire  _GEN_366 = 3'h3 == _rs2ROBEntry_T_7[2:0] ? io_robRead_3_busy : _GEN_365; // @[ReservationStation.scala 181:{48,48}]
  wire  _GEN_367 = 3'h4 == _rs2ROBEntry_T_7[2:0] ? io_robRead_4_busy : _GEN_366; // @[ReservationStation.scala 181:{48,48}]
  wire [4:0] _GEN_369 = 3'h1 == _rs2ROBEntry_T_7[2:0] ? io_robRead_1_rd : io_robRead_0_rd; // @[ReservationStation.scala 181:{132,132}]
  wire [4:0] _GEN_370 = 3'h2 == _rs2ROBEntry_T_7[2:0] ? io_robRead_2_rd : _GEN_369; // @[ReservationStation.scala 181:{132,132}]
  wire [4:0] _GEN_371 = 3'h3 == _rs2ROBEntry_T_7[2:0] ? io_robRead_3_rd : _GEN_370; // @[ReservationStation.scala 181:{132,132}]
  wire [4:0] _GEN_372 = 3'h4 == _rs2ROBEntry_T_7[2:0] ? io_robRead_4_rd : _GEN_371; // @[ReservationStation.scala 181:{132,132}]
  wire  rs2FromROB_2 = (_GEN_367 & _GEN_362 == 2'h2 | _GEN_362 == 2'h3) & _GEN_372 == entries_2_rs2 & entries_2_rs2 != 5'h0
    ; // @[ReservationStation.scala 181:142]
  wire  _T_24 = entries_2_rs1ROBId != 8'h0; // @[ReservationStation.scala 182:43]
  wire [31:0] _GEN_374 = 3'h1 == _rs1ROBEntry_T_7[2:0] ? io_robRead_1_data : io_robRead_0_data; // @[ReservationStation.scala 183:{26,26}]
  wire [31:0] _GEN_375 = 3'h2 == _rs1ROBEntry_T_7[2:0] ? io_robRead_2_data : _GEN_374; // @[ReservationStation.scala 183:{26,26}]
  wire [31:0] _GEN_376 = 3'h3 == _rs1ROBEntry_T_7[2:0] ? io_robRead_3_data : _GEN_375; // @[ReservationStation.scala 183:{26,26}]
  wire  _T_26 = entries_2_rs2ROBId != 8'h0; // @[ReservationStation.scala 186:43]
  wire [31:0] _GEN_381 = 3'h1 == _rs2ROBEntry_T_7[2:0] ? io_robRead_1_data : io_robRead_0_data; // @[ReservationStation.scala 187:{26,26}]
  wire [31:0] _GEN_382 = 3'h2 == _rs2ROBEntry_T_7[2:0] ? io_robRead_2_data : _GEN_381; // @[ReservationStation.scala 187:{26,26}]
  wire [31:0] _GEN_383 = 3'h3 == _rs2ROBEntry_T_7[2:0] ? io_robRead_3_data : _GEN_382; // @[ReservationStation.scala 187:{26,26}]
  wire  _rs1MatchVec_T_8 = io_cdb_0_bits_rd == entries_2_rs1; // @[ReservationStation.scala 192:61]
  wire  _rs1MatchVec_T_9 = io_cdb_1_bits_rd == entries_2_rs1; // @[ReservationStation.scala 192:61]
  wire  _rs1MatchVec_T_10 = io_cdb_2_bits_rd == entries_2_rs1; // @[ReservationStation.scala 192:61]
  wire  _rs1MatchVec_T_11 = io_cdb_3_bits_rd == entries_2_rs1; // @[ReservationStation.scala 192:61]
  wire [3:0] rs1MatchVec_2 = {_rs1MatchVec_T_11,_rs1MatchVec_T_10,_rs1MatchVec_T_9,_rs1MatchVec_T_8}; // @[Cat.scala 33:92]
  wire  _rs2MatchVec_T_8 = io_cdb_0_bits_rd == entries_2_rs2; // @[ReservationStation.scala 193:61]
  wire  _rs2MatchVec_T_9 = io_cdb_1_bits_rd == entries_2_rs2; // @[ReservationStation.scala 193:61]
  wire  _rs2MatchVec_T_10 = io_cdb_2_bits_rd == entries_2_rs2; // @[ReservationStation.scala 193:61]
  wire  _rs2MatchVec_T_11 = io_cdb_3_bits_rd == entries_2_rs2; // @[ReservationStation.scala 193:61]
  wire [3:0] rs2MatchVec_2 = {_rs2MatchVec_T_11,_rs2MatchVec_T_10,_rs2MatchVec_T_9,_rs2MatchVec_T_8}; // @[Cat.scala 33:92]
  wire  _rs1IDMatchVec_T_8 = io_cdb_0_bits_id == entries_2_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire  _rs1IDMatchVec_T_9 = io_cdb_1_bits_id == entries_2_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire  _rs1IDMatchVec_T_10 = io_cdb_2_bits_id == entries_2_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire  _rs1IDMatchVec_T_11 = io_cdb_3_bits_id == entries_2_rs1ROBId; // @[ReservationStation.scala 194:63]
  wire [3:0] rs1IDMatchVec_2 = {_rs1IDMatchVec_T_11,_rs1IDMatchVec_T_10,_rs1IDMatchVec_T_9,_rs1IDMatchVec_T_8}; // @[Cat.scala 33:92]
  wire  _rs2IDMatchVec_T_8 = io_cdb_0_bits_id == entries_2_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire  _rs2IDMatchVec_T_9 = io_cdb_1_bits_id == entries_2_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire  _rs2IDMatchVec_T_10 = io_cdb_2_bits_id == entries_2_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire  _rs2IDMatchVec_T_11 = io_cdb_3_bits_id == entries_2_rs2ROBId; // @[ReservationStation.scala 195:63]
  wire [3:0] rs2IDMatchVec_2 = {_rs2IDMatchVec_T_11,_rs2IDMatchVec_T_10,_rs2IDMatchVec_T_9,_rs2IDMatchVec_T_8}; // @[Cat.scala 33:92]
  wire [3:0] _cdbBypassRs1_T_2 = cdbValidVec & rs1MatchVec_2; // @[ReservationStation.scala 197:44]
  wire [3:0] cdbBypassRs1_2 = _cdbBypassRs1_T_2 & rs1IDMatchVec_2; // @[ReservationStation.scala 197:58]
  wire [3:0] _cdbBypassRs2_T_2 = cdbValidVec & rs2MatchVec_2; // @[ReservationStation.scala 198:44]
  wire [3:0] cdbBypassRs2_2 = _cdbBypassRs2_T_2 & rs2IDMatchVec_2; // @[ReservationStation.scala 198:58]
  wire  bypassRs1_2 = |cdbBypassRs1_2; // @[ReservationStation.scala 200:42]
  wire  bypassRs2_2 = |cdbBypassRs2_2; // @[ReservationStation.scala 201:42]
  wire [31:0] _entries_2_rs1Val_T_4 = cdbBypassRs1_2[0] ? io_cdb_0_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs1Val_T_5 = cdbBypassRs1_2[1] ? io_cdb_1_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs1Val_T_6 = cdbBypassRs1_2[2] ? io_cdb_2_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs1Val_T_7 = cdbBypassRs1_2[3] ? io_cdb_3_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs1Val_T_8 = _entries_2_rs1Val_T_4 | _entries_2_rs1Val_T_5; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs1Val_T_9 = _entries_2_rs1Val_T_8 | _entries_2_rs1Val_T_6; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs1Val_T_10 = _entries_2_rs1Val_T_9 | _entries_2_rs1Val_T_7; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs2Val_T_4 = cdbBypassRs2_2[0] ? io_cdb_0_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs2Val_T_5 = cdbBypassRs2_2[1] ? io_cdb_1_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs2Val_T_6 = cdbBypassRs2_2[2] ? io_cdb_2_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs2Val_T_7 = cdbBypassRs2_2[3] ? io_cdb_3_bits_data : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs2Val_T_8 = _entries_2_rs2Val_T_4 | _entries_2_rs2Val_T_5; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs2Val_T_9 = _entries_2_rs2Val_T_8 | _entries_2_rs2Val_T_6; // @[Mux.scala 27:73]
  wire [31:0] _entries_2_rs2Val_T_10 = _entries_2_rs2Val_T_9 | _entries_2_rs2Val_T_7; // @[Mux.scala 27:73]
  assign io_enq_ready = ~full & ~_GEN_8; // @[ReservationStation.scala 95:27]
  assign io_deq_valid = oprReady & _GEN_11; // @[ReservationStation.scala 96:30]
  assign io_deq_bits_op = 2'h2 == head ? entries_2_op : _GEN_13; // @[ReservationStation.scala 97:{20,20}]
  assign io_deq_bits_ROBId = 2'h2 == head ? entries_2_ROBId : _GEN_16; // @[ReservationStation.scala 98:{23,23}]
  assign io_deq_bits_opr1 = 2'h2 == head ? entries_2_opr1 : _GEN_19; // @[ReservationStation.scala 99:{22,22}]
  assign io_deq_bits_opr2 = 2'h2 == head ? entries_2_opr2 : _GEN_22; // @[ReservationStation.scala 100:{22,22}]
  assign io_deq_bits_rs1Val = 2'h2 == head ? entries_2_rs1Val : _GEN_25; // @[ReservationStation.scala 101:{24,24}]
  assign io_deq_bits_rs2Val = 2'h2 == head ? entries_2_rs2Val : _GEN_28; // @[ReservationStation.scala 102:{24,24}]
  assign io_deq_bits_immSrc = 2'h2 == head ? entries_2_immSrc : _GEN_31; // @[ReservationStation.scala 103:{24,24}]
  assign io_deq_bits_immSign = 2'h2 == head ? entries_2_immSign : _GEN_34; // @[ReservationStation.scala 104:{25,25}]
  assign io_deq_bits_excpType = 2'h2 == head ? entries_2_excpType : _GEN_37; // @[ReservationStation.scala 105:{26,26}]
  assign io_deq_bits_pc = 2'h2 == head ? entries_2_pc : _GEN_40; // @[ReservationStation.scala 106:{20,20}]
  assign io_deq_bits_inst = 2'h2 == head ? entries_2_inst : _GEN_43; // @[ReservationStation.scala 107:{22,22}]
  assign io_robOut_valid = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign io_robOut_bits_id = _GEN_233[2:0];
  assign io_rf_0_addr = _T ? io_enq_bits_rs1 : 5'h0; // @[ReservationStation.scala 115:16 120:24 144:23]
  assign io_rf_1_addr = _T ? io_enq_bits_rs2 : 5'h0; // @[ReservationStation.scala 115:16 120:24 145:23]
  always @(posedge clock) begin
    if (io_flush) begin // @[ReservationStation.scala 213:21]
      entries_0_busy <= 1'h0; // @[ReservationStation.scala 214:37]
    end else if (_T_1) begin // @[ReservationStation.scala 152:24]
      if (2'h0 == head) begin // @[ReservationStation.scala 153:28]
        entries_0_busy <= 1'h0; // @[ReservationStation.scala 153:28]
      end else begin
        entries_0_busy <= _GEN_169;
      end
    end else begin
      entries_0_busy <= _GEN_169;
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 123:26]
        entries_0_op <= io_enq_bits_op; // @[ReservationStation.scala 123:26]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 122:29]
        entries_0_ROBId <= io_enq_bits_ROBId; // @[ReservationStation.scala 122:29]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 127:28]
        entries_0_opr1 <= io_enq_bits_opr1; // @[ReservationStation.scala 127:28]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 128:28]
        entries_0_opr2 <= io_enq_bits_opr2; // @[ReservationStation.scala 128:28]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 129:27]
        entries_0_rs1 <= io_enq_bits_rs1; // @[ReservationStation.scala 129:27]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 130:27]
        entries_0_rs2 <= io_enq_bits_rs2; // @[ReservationStation.scala 130:27]
      end
    end
    if (entries_0_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs1 & _T_8) begin // @[ReservationStation.scala 202:51]
        entries_0_rs1Val <= _entries_0_rs1Val_T_10; // @[ReservationStation.scala 203:26]
      end else if (rs1FromROB & entries_0_rs1ROBId != 8'h0) begin // @[ReservationStation.scala 182:52]
        if (3'h4 == _rs1ROBEntry_T_1[2:0]) begin // @[ReservationStation.scala 183:26]
          entries_0_rs1Val <= io_robRead_4_data; // @[ReservationStation.scala 183:26]
        end else begin
          entries_0_rs1Val <= _GEN_272;
        end
      end else begin
        entries_0_rs1Val <= _GEN_216;
      end
    end else begin
      entries_0_rs1Val <= _GEN_216;
    end
    if (entries_0_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs2 & _T_10) begin // @[ReservationStation.scala 206:51]
        entries_0_rs2Val <= _entries_0_rs2Val_T_10; // @[ReservationStation.scala 207:26]
      end else if (rs2FromROB & entries_0_rs2ROBId != 8'h0) begin // @[ReservationStation.scala 186:52]
        if (3'h4 == _rs2ROBEntry_T_1[2:0]) begin // @[ReservationStation.scala 187:26]
          entries_0_rs2Val <= io_robRead_4_data; // @[ReservationStation.scala 187:26]
        end else begin
          entries_0_rs2Val <= _GEN_279;
        end
      end else begin
        entries_0_rs2Val <= _GEN_219;
      end
    end else begin
      entries_0_rs2Val <= _GEN_219;
    end
    if (entries_0_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs1 & _T_8) begin // @[ReservationStation.scala 202:51]
        entries_0_rs1ROBId <= 8'h0; // @[ReservationStation.scala 204:28]
      end else if (rs1FromROB & entries_0_rs1ROBId != 8'h0) begin // @[ReservationStation.scala 182:52]
        entries_0_rs1ROBId <= 8'h0; // @[ReservationStation.scala 184:28]
      end else begin
        entries_0_rs1ROBId <= _GEN_178;
      end
    end else begin
      entries_0_rs1ROBId <= _GEN_178;
    end
    if (entries_0_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs2 & _T_10) begin // @[ReservationStation.scala 206:51]
        entries_0_rs2ROBId <= 8'h0; // @[ReservationStation.scala 208:28]
      end else if (rs2FromROB & entries_0_rs2ROBId != 8'h0) begin // @[ReservationStation.scala 186:52]
        entries_0_rs2ROBId <= 8'h0; // @[ReservationStation.scala 188:28]
      end else begin
        entries_0_rs2ROBId <= _GEN_181;
      end
    end else begin
      entries_0_rs2ROBId <= _GEN_181;
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 132:30]
        entries_0_immSrc <= io_enq_bits_immSrc; // @[ReservationStation.scala 132:30]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 133:31]
        entries_0_immSign <= io_enq_bits_immSign; // @[ReservationStation.scala 133:31]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 134:32]
        entries_0_excpType <= io_enq_bits_excpType; // @[ReservationStation.scala 134:32]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 135:26]
        entries_0_pc <= io_enq_bits_pc; // @[ReservationStation.scala 135:26]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h0 == tail) begin // @[ReservationStation.scala 136:28]
        entries_0_inst <= io_enq_bits_inst; // @[ReservationStation.scala 136:28]
      end else if (2'h0 == tail) begin // @[ReservationStation.scala 126:28]
        entries_0_inst <= io_enq_bits_inst; // @[ReservationStation.scala 126:28]
      end
    end
    if (io_flush) begin // @[ReservationStation.scala 213:21]
      entries_1_busy <= 1'h0; // @[ReservationStation.scala 214:37]
    end else if (_T_1) begin // @[ReservationStation.scala 152:24]
      if (2'h1 == head) begin // @[ReservationStation.scala 153:28]
        entries_1_busy <= 1'h0; // @[ReservationStation.scala 153:28]
      end else begin
        entries_1_busy <= _GEN_170;
      end
    end else begin
      entries_1_busy <= _GEN_170;
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 123:26]
        entries_1_op <= io_enq_bits_op; // @[ReservationStation.scala 123:26]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 122:29]
        entries_1_ROBId <= io_enq_bits_ROBId; // @[ReservationStation.scala 122:29]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 127:28]
        entries_1_opr1 <= io_enq_bits_opr1; // @[ReservationStation.scala 127:28]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 128:28]
        entries_1_opr2 <= io_enq_bits_opr2; // @[ReservationStation.scala 128:28]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 129:27]
        entries_1_rs1 <= io_enq_bits_rs1; // @[ReservationStation.scala 129:27]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 130:27]
        entries_1_rs2 <= io_enq_bits_rs2; // @[ReservationStation.scala 130:27]
      end
    end
    if (entries_1_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs1_1 & _T_16) begin // @[ReservationStation.scala 202:51]
        entries_1_rs1Val <= _entries_1_rs1Val_T_10; // @[ReservationStation.scala 203:26]
      end else if (rs1FromROB_1 & entries_1_rs1ROBId != 8'h0) begin // @[ReservationStation.scala 182:52]
        if (3'h4 == _rs1ROBEntry_T_4[2:0]) begin // @[ReservationStation.scala 183:26]
          entries_1_rs1Val <= io_robRead_4_data; // @[ReservationStation.scala 183:26]
        end else begin
          entries_1_rs1Val <= _GEN_324;
        end
      end else begin
        entries_1_rs1Val <= _GEN_217;
      end
    end else begin
      entries_1_rs1Val <= _GEN_217;
    end
    if (entries_1_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs2_1 & _T_18) begin // @[ReservationStation.scala 206:51]
        entries_1_rs2Val <= _entries_1_rs2Val_T_10; // @[ReservationStation.scala 207:26]
      end else if (rs2FromROB_1 & entries_1_rs2ROBId != 8'h0) begin // @[ReservationStation.scala 186:52]
        if (3'h4 == _rs2ROBEntry_T_4[2:0]) begin // @[ReservationStation.scala 187:26]
          entries_1_rs2Val <= io_robRead_4_data; // @[ReservationStation.scala 187:26]
        end else begin
          entries_1_rs2Val <= _GEN_331;
        end
      end else begin
        entries_1_rs2Val <= _GEN_220;
      end
    end else begin
      entries_1_rs2Val <= _GEN_220;
    end
    if (entries_1_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs1_1 & _T_16) begin // @[ReservationStation.scala 202:51]
        entries_1_rs1ROBId <= 8'h0; // @[ReservationStation.scala 204:28]
      end else if (rs1FromROB_1 & entries_1_rs1ROBId != 8'h0) begin // @[ReservationStation.scala 182:52]
        entries_1_rs1ROBId <= 8'h0; // @[ReservationStation.scala 184:28]
      end else begin
        entries_1_rs1ROBId <= _GEN_179;
      end
    end else begin
      entries_1_rs1ROBId <= _GEN_179;
    end
    if (entries_1_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs2_1 & _T_18) begin // @[ReservationStation.scala 206:51]
        entries_1_rs2ROBId <= 8'h0; // @[ReservationStation.scala 208:28]
      end else if (rs2FromROB_1 & entries_1_rs2ROBId != 8'h0) begin // @[ReservationStation.scala 186:52]
        entries_1_rs2ROBId <= 8'h0; // @[ReservationStation.scala 188:28]
      end else begin
        entries_1_rs2ROBId <= _GEN_182;
      end
    end else begin
      entries_1_rs2ROBId <= _GEN_182;
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 132:30]
        entries_1_immSrc <= io_enq_bits_immSrc; // @[ReservationStation.scala 132:30]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 133:31]
        entries_1_immSign <= io_enq_bits_immSign; // @[ReservationStation.scala 133:31]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 134:32]
        entries_1_excpType <= io_enq_bits_excpType; // @[ReservationStation.scala 134:32]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 135:26]
        entries_1_pc <= io_enq_bits_pc; // @[ReservationStation.scala 135:26]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h1 == tail) begin // @[ReservationStation.scala 136:28]
        entries_1_inst <= io_enq_bits_inst; // @[ReservationStation.scala 136:28]
      end else if (2'h1 == tail) begin // @[ReservationStation.scala 126:28]
        entries_1_inst <= io_enq_bits_inst; // @[ReservationStation.scala 126:28]
      end
    end
    if (io_flush) begin // @[ReservationStation.scala 213:21]
      entries_2_busy <= 1'h0; // @[ReservationStation.scala 214:37]
    end else if (_T_1) begin // @[ReservationStation.scala 152:24]
      if (2'h2 == head) begin // @[ReservationStation.scala 153:28]
        entries_2_busy <= 1'h0; // @[ReservationStation.scala 153:28]
      end else begin
        entries_2_busy <= _GEN_171;
      end
    end else begin
      entries_2_busy <= _GEN_171;
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 123:26]
        entries_2_op <= io_enq_bits_op; // @[ReservationStation.scala 123:26]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 122:29]
        entries_2_ROBId <= io_enq_bits_ROBId; // @[ReservationStation.scala 122:29]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 127:28]
        entries_2_opr1 <= io_enq_bits_opr1; // @[ReservationStation.scala 127:28]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 128:28]
        entries_2_opr2 <= io_enq_bits_opr2; // @[ReservationStation.scala 128:28]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 129:27]
        entries_2_rs1 <= io_enq_bits_rs1; // @[ReservationStation.scala 129:27]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 130:27]
        entries_2_rs2 <= io_enq_bits_rs2; // @[ReservationStation.scala 130:27]
      end
    end
    if (entries_2_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs1_2 & _T_24) begin // @[ReservationStation.scala 202:51]
        entries_2_rs1Val <= _entries_2_rs1Val_T_10; // @[ReservationStation.scala 203:26]
      end else if (rs1FromROB_2 & entries_2_rs1ROBId != 8'h0) begin // @[ReservationStation.scala 182:52]
        if (3'h4 == _rs1ROBEntry_T_7[2:0]) begin // @[ReservationStation.scala 183:26]
          entries_2_rs1Val <= io_robRead_4_data; // @[ReservationStation.scala 183:26]
        end else begin
          entries_2_rs1Val <= _GEN_376;
        end
      end else begin
        entries_2_rs1Val <= _GEN_218;
      end
    end else begin
      entries_2_rs1Val <= _GEN_218;
    end
    if (entries_2_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs2_2 & _T_26) begin // @[ReservationStation.scala 206:51]
        entries_2_rs2Val <= _entries_2_rs2Val_T_10; // @[ReservationStation.scala 207:26]
      end else if (rs2FromROB_2 & entries_2_rs2ROBId != 8'h0) begin // @[ReservationStation.scala 186:52]
        if (3'h4 == _rs2ROBEntry_T_7[2:0]) begin // @[ReservationStation.scala 187:26]
          entries_2_rs2Val <= io_robRead_4_data; // @[ReservationStation.scala 187:26]
        end else begin
          entries_2_rs2Val <= _GEN_383;
        end
      end else begin
        entries_2_rs2Val <= _GEN_221;
      end
    end else begin
      entries_2_rs2Val <= _GEN_221;
    end
    if (entries_2_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs1_2 & _T_24) begin // @[ReservationStation.scala 202:51]
        entries_2_rs1ROBId <= 8'h0; // @[ReservationStation.scala 204:28]
      end else if (rs1FromROB_2 & entries_2_rs1ROBId != 8'h0) begin // @[ReservationStation.scala 182:52]
        entries_2_rs1ROBId <= 8'h0; // @[ReservationStation.scala 184:28]
      end else begin
        entries_2_rs1ROBId <= _GEN_180;
      end
    end else begin
      entries_2_rs1ROBId <= _GEN_180;
    end
    if (entries_2_busy) begin // @[ReservationStation.scala 171:22]
      if (bypassRs2_2 & _T_26) begin // @[ReservationStation.scala 206:51]
        entries_2_rs2ROBId <= 8'h0; // @[ReservationStation.scala 208:28]
      end else if (rs2FromROB_2 & entries_2_rs2ROBId != 8'h0) begin // @[ReservationStation.scala 186:52]
        entries_2_rs2ROBId <= 8'h0; // @[ReservationStation.scala 188:28]
      end else begin
        entries_2_rs2ROBId <= _GEN_183;
      end
    end else begin
      entries_2_rs2ROBId <= _GEN_183;
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 132:30]
        entries_2_immSrc <= io_enq_bits_immSrc; // @[ReservationStation.scala 132:30]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 133:31]
        entries_2_immSign <= io_enq_bits_immSign; // @[ReservationStation.scala 133:31]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 134:32]
        entries_2_excpType <= io_enq_bits_excpType; // @[ReservationStation.scala 134:32]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 135:26]
        entries_2_pc <= io_enq_bits_pc; // @[ReservationStation.scala 135:26]
      end
    end
    if (_T) begin // @[ReservationStation.scala 120:24]
      if (2'h2 == tail) begin // @[ReservationStation.scala 136:28]
        entries_2_inst <= io_enq_bits_inst; // @[ReservationStation.scala 136:28]
      end else if (2'h2 == tail) begin // @[ReservationStation.scala 126:28]
        entries_2_inst <= io_enq_bits_inst; // @[ReservationStation.scala 126:28]
      end
    end
    if (reset) begin // @[ReservationStation.scala 86:23]
      head <= 2'h0; // @[ReservationStation.scala 86:23]
    end else if (io_flush) begin // @[ReservationStation.scala 213:21]
      head <= 2'h0; // @[ReservationStation.scala 215:14]
    end else if (_T_1) begin // @[ReservationStation.scala 152:24]
      if (head == 2'h2) begin // @[ReservationStation.scala 158:20]
        head <= 2'h0;
      end else begin
        head <= _head_T_2;
      end
    end
    if (reset) begin // @[ReservationStation.scala 87:23]
      tail <= 2'h0; // @[ReservationStation.scala 87:23]
    end else if (io_flush) begin // @[ReservationStation.scala 213:21]
      tail <= 2'h0; // @[ReservationStation.scala 216:14]
    end else if (_T) begin // @[ReservationStation.scala 120:24]
      if (tail == 2'h2) begin // @[ReservationStation.scala 149:20]
        tail <= 2'h0;
      end else begin
        tail <= _tail_T_2;
      end
    end
    if (reset) begin // @[ReservationStation.scala 89:24]
      count <= 2'h0; // @[ReservationStation.scala 89:24]
    end else if (io_flush) begin // @[ReservationStation.scala 213:21]
      count <= 2'h0; // @[ReservationStation.scala 217:15]
    end else if (~(_T_1 & _T)) begin // @[ReservationStation.scala 161:43]
      if (_T_1) begin // @[ReservationStation.scala 165:27]
        count <= _count_T_3; // @[ReservationStation.scala 166:19]
      end else begin
        count <= _GEN_236;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  entries_0_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  entries_0_op = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  entries_0_ROBId = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  entries_0_opr1 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  entries_0_opr2 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  entries_0_rs1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  entries_0_rs2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  entries_0_rs1Val = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  entries_0_rs2Val = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  entries_0_rs1ROBId = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  entries_0_rs2ROBId = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  entries_0_immSrc = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  entries_0_immSign = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  entries_0_excpType = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  entries_0_pc = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  entries_0_inst = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  entries_1_busy = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  entries_1_op = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  entries_1_ROBId = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  entries_1_opr1 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  entries_1_opr2 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  entries_1_rs1 = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  entries_1_rs2 = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  entries_1_rs1Val = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  entries_1_rs2Val = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  entries_1_rs1ROBId = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  entries_1_rs2ROBId = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  entries_1_immSrc = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  entries_1_immSign = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  entries_1_excpType = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  entries_1_pc = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  entries_1_inst = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  entries_2_busy = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  entries_2_op = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  entries_2_ROBId = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  entries_2_opr1 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  entries_2_opr2 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  entries_2_rs1 = _RAND_37[4:0];
  _RAND_38 = {1{`RANDOM}};
  entries_2_rs2 = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  entries_2_rs1Val = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  entries_2_rs2Val = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  entries_2_rs1ROBId = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  entries_2_rs2ROBId = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  entries_2_immSrc = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  entries_2_immSign = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  entries_2_excpType = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  entries_2_pc = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  entries_2_inst = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  head = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  tail = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  count = _RAND_50[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BRU(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  input  [31:0] io_offset,
  input  [31:0] io_pc,
  input  [3:0]  io_opSel,
  output [31:0] io_brAddr,
  output        io_brTaken
);
  wire  _cmp_T_2 = $signed(io_in1) < $signed(io_in2); // @[BRU.scala 30:47]
  wire  _cmp_T_3 = io_in1 < io_in2; // @[BRU.scala 31:40]
  wire  _cmp_T_4 = io_in1 == io_in2; // @[BRU.scala 32:40]
  wire  _cmp_T_5 = io_in1 != io_in2; // @[BRU.scala 33:40]
  wire  _cmp_T_8 = $signed(io_in1) >= $signed(io_in2); // @[BRU.scala 34:47]
  wire  _cmp_T_9 = io_in1 >= io_in2; // @[BRU.scala 35:40]
  wire  _cmp_T_13 = 4'h7 == io_opSel ? _cmp_T_3 : 4'h6 == io_opSel & _cmp_T_2; // @[Mux.scala 81:58]
  wire  _cmp_T_15 = 4'h3 == io_opSel ? _cmp_T_4 : _cmp_T_13; // @[Mux.scala 81:58]
  wire  _cmp_T_17 = 4'h4 == io_opSel ? _cmp_T_5 : _cmp_T_15; // @[Mux.scala 81:58]
  wire  _cmp_T_19 = 4'h5 == io_opSel ? _cmp_T_8 : _cmp_T_17; // @[Mux.scala 81:58]
  wire  cmp = 4'h8 == io_opSel ? _cmp_T_9 : _cmp_T_19; // @[Mux.scala 81:58]
  wire  _T = io_opSel == 4'h1; // @[BRU.scala 39:19]
  wire [31:0] _brAddr_T_1 = io_pc + io_offset; // @[BRU.scala 40:25]
  wire  _T_1 = io_opSel == 4'h2; // @[BRU.scala 41:25]
  wire [31:0] _brAddr_T_3 = io_in1 + io_offset; // @[BRU.scala 42:26]
  wire [31:0] _GEN_0 = cmp ? _brAddr_T_1 : _brAddr_T_1; // @[BRU.scala 43:32 44:16 46:16]
  wire [31:0] _GEN_1 = io_opSel == 4'h2 ? _brAddr_T_3 : _GEN_0; // @[BRU.scala 41:38 42:16]
  assign io_brAddr = io_opSel == 4'h1 ? _brAddr_T_1 : _GEN_1; // @[BRU.scala 39:31 40:16]
  assign io_brTaken = cmp | _T | _T_1; // @[BRU.scala 50:45]
endmodule
module BRUStage_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [3:0]  io_in_bits_opr1,
  input  [3:0]  io_in_bits_opr2,
  input  [3:0]  io_in_bits_bruOp,
  input  [2:0]  io_in_bits_immSrc,
  input  [31:0] io_in_bits_rs1Val,
  input  [31:0] io_in_bits_rs2Val,
  input  [31:0] io_in_bits_inst,
  input  [31:0] io_in_bits_pc,
  input  [7:0]  io_in_bits_id,
  output        io_out_valid,
  output        io_out_bits_brTaken,
  output [31:0] io_out_bits_brAddr,
  output [4:0]  io_out_bits_rd,
  output [31:0] io_out_bits_data,
  output [7:0]  io_out_bits_id,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] immGen_io_inst; // @[BRU.scala 228:24]
  wire [2:0] immGen_io_immSrc; // @[BRU.scala 228:24]
  wire  immGen_io_immSign; // @[BRU.scala 228:24]
  wire [31:0] immGen_io_imm; // @[BRU.scala 228:24]
  wire [31:0] bru_io_in1; // @[BRU.scala 263:21]
  wire [31:0] bru_io_in2; // @[BRU.scala 263:21]
  wire [31:0] bru_io_offset; // @[BRU.scala 263:21]
  wire [31:0] bru_io_pc; // @[BRU.scala 263:21]
  wire [3:0] bru_io_opSel; // @[BRU.scala 263:21]
  wire [31:0] bru_io_brAddr; // @[BRU.scala 263:21]
  wire  bru_io_brTaken; // @[BRU.scala 263:21]
  reg  s0_full; // @[BRU.scala 220:26]
  reg  s1_full; // @[BRU.scala 250:26]
  wire  s1_ready = ~s1_full | io_out_valid; // @[BRU.scala 258:26]
  wire  s0_fire = s0_full & s1_ready; // @[BRU.scala 221:28]
  wire  s0_ready = ~s0_full | s0_fire; // @[BRU.scala 223:26]
  wire  s0_latch = io_in_valid & s0_ready; // @[BRU.scala 219:32]
  reg [3:0] s0_info_opr1; // @[Reg.scala 19:16]
  reg [3:0] s0_info_opr2; // @[Reg.scala 19:16]
  reg [3:0] s0_info_bruOp; // @[Reg.scala 19:16]
  reg [2:0] s0_info_immSrc; // @[Reg.scala 19:16]
  reg [31:0] s0_info_rs1Val; // @[Reg.scala 19:16]
  reg [31:0] s0_info_rs2Val; // @[Reg.scala 19:16]
  reg [31:0] s0_info_inst; // @[Reg.scala 19:16]
  reg [31:0] s0_info_pc; // @[Reg.scala 19:16]
  reg [7:0] s0_info_id; // @[Reg.scala 19:16]
  wire  _GEN_9 = s0_fire & s0_full ? 1'h0 : s0_full; // @[BRU.scala 220:26 226:{35,45}]
  wire  _GEN_10 = s0_latch | _GEN_9; // @[BRU.scala 225:{20,30}]
  reg [3:0] s1_bruOp; // @[Reg.scala 19:16]
  reg [31:0] s1_bruInVec_0; // @[Reg.scala 19:16]
  reg [31:0] s1_bruInVec_1; // @[Reg.scala 19:16]
  reg [31:0] s1_imm; // @[Reg.scala 19:16]
  reg [31:0] s1_pc; // @[Reg.scala 19:16]
  reg [31:0] s1_inst; // @[Reg.scala 19:16]
  reg [7:0] s1_id; // @[Reg.scala 19:16]
  wire  _GEN_18 = io_out_valid & s1_full ? 1'h0 : s1_full; // @[BRU.scala 250:26 261:{35,45}]
  wire  _GEN_19 = s0_fire | _GEN_18; // @[BRU.scala 260:{20,30}]
  ImmGen immGen ( // @[BRU.scala 228:24]
    .io_inst(immGen_io_inst),
    .io_immSrc(immGen_io_immSrc),
    .io_immSign(immGen_io_immSign),
    .io_imm(immGen_io_imm)
  );
  BRU bru ( // @[BRU.scala 263:21]
    .io_in1(bru_io_in1),
    .io_in2(bru_io_in2),
    .io_offset(bru_io_offset),
    .io_pc(bru_io_pc),
    .io_opSel(bru_io_opSel),
    .io_brAddr(bru_io_brAddr),
    .io_brTaken(bru_io_brTaken)
  );
  assign io_in_ready = ~s0_full | s0_fire; // @[BRU.scala 223:26]
  assign io_out_valid = s1_full; // @[BRU.scala 276:18]
  assign io_out_bits_brTaken = bru_io_brTaken & s1_full; // @[BRU.scala 270:43]
  assign io_out_bits_brAddr = bru_io_brAddr; // @[BRU.scala 271:24]
  assign io_out_bits_rd = s1_bruOp != 4'h2 | s1_bruOp != 4'h1 ? 5'h0 : s1_inst[11:7]; // @[BRU.scala 272:26]
  assign io_out_bits_data = s1_pc + 32'h4; // @[BRU.scala 274:31]
  assign io_out_bits_id = s1_id; // @[BRU.scala 275:20]
  assign immGen_io_inst = s0_info_inst; // @[BRU.scala 232:20]
  assign immGen_io_immSrc = s0_info_immSrc; // @[BRU.scala 230:22]
  assign immGen_io_immSign = 1'h1; // @[BRU.scala 231:23]
  assign bru_io_in1 = s1_bruInVec_0; // @[BRU.scala 264:16]
  assign bru_io_in2 = s1_bruInVec_1; // @[BRU.scala 265:16]
  assign bru_io_offset = s1_imm; // @[BRU.scala 266:19]
  assign bru_io_pc = s1_pc; // @[BRU.scala 267:15]
  assign bru_io_opSel = s1_bruOp; // @[BRU.scala 268:18]
  always @(posedge clock) begin
    if (reset) begin // @[BRU.scala 220:26]
      s0_full <= 1'h0; // @[BRU.scala 220:26]
    end else if (io_flush) begin // @[BRU.scala 280:20]
      s0_full <= 1'h0; // @[BRU.scala 281:17]
    end else begin
      s0_full <= _GEN_10;
    end
    if (reset) begin // @[BRU.scala 250:26]
      s1_full <= 1'h0; // @[BRU.scala 250:26]
    end else if (io_flush) begin // @[BRU.scala 280:20]
      s1_full <= 1'h0; // @[BRU.scala 282:17]
    end else begin
      s1_full <= _GEN_19;
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_opr1 <= io_in_bits_opr1; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_opr2 <= io_in_bits_opr2; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_bruOp <= io_in_bits_bruOp; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_immSrc <= io_in_bits_immSrc; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_rs1Val <= io_in_bits_rs1Val; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_rs2Val <= io_in_bits_rs2Val; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_inst <= io_in_bits_inst; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_pc <= io_in_bits_pc; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_id <= io_in_bits_id; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_bruOp <= s0_info_bruOp; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      if (4'h1 == s0_info_opr1) begin // @[Mux.scala 81:58]
        s1_bruInVec_0 <= s0_info_rs1Val;
      end else begin
        s1_bruInVec_0 <= 32'h0;
      end
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      if (4'h2 == s0_info_opr2) begin // @[Mux.scala 81:58]
        s1_bruInVec_1 <= s0_info_rs2Val;
      end else begin
        s1_bruInVec_1 <= 32'h0;
      end
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_imm <= immGen_io_imm; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_pc <= s0_info_pc; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_inst <= s0_info_inst; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_id <= s0_info_id; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s1_full = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s0_info_opr1 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  s0_info_opr2 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  s0_info_bruOp = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  s0_info_immSrc = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  s0_info_rs1Val = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  s0_info_rs2Val = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  s0_info_inst = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  s0_info_pc = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  s0_info_id = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  s1_bruOp = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  s1_bruInVec_0 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  s1_bruInVec_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  s1_imm = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  s1_pc = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  s1_inst = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  s1_id = _RAND_17[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSUQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_decInfo_en,
  input         io_enq_bits_decInfo_wen,
  input         io_enq_bits_decInfo_load,
  input  [1:0]  io_enq_bits_decInfo_wd,
  input         io_enq_bits_decInfo_signed,
  input  [31:0] io_enq_bits_addr,
  input  [31:0] io_enq_bits_rs2Val,
  input  [7:0]  io_enq_bits_id,
  input  [4:0]  io_enq_bits_rd,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_decInfo_en,
  output        io_deq_bits_decInfo_wen,
  output        io_deq_bits_decInfo_load,
  output [1:0]  io_deq_bits_decInfo_wd,
  output        io_deq_bits_decInfo_signed,
  output [31:0] io_deq_bits_addr,
  output [31:0] io_deq_bits_rs2Val,
  output [7:0]  io_deq_bits_id,
  output [4:0]  io_deq_bits_rd,
  input  [7:0]  io_rob_bits_id,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
`endif // RANDOMIZE_REG_INIT
  reg  entries_0_busy; // @[LSUQueue.scala 43:22]
  reg  entries_0_ready; // @[LSUQueue.scala 43:22]
  reg  entries_0_decInfo_en; // @[LSUQueue.scala 43:22]
  reg  entries_0_decInfo_wen; // @[LSUQueue.scala 43:22]
  reg  entries_0_decInfo_load; // @[LSUQueue.scala 43:22]
  reg [1:0] entries_0_decInfo_wd; // @[LSUQueue.scala 43:22]
  reg  entries_0_decInfo_signed; // @[LSUQueue.scala 43:22]
  reg [31:0] entries_0_addr; // @[LSUQueue.scala 43:22]
  reg [31:0] entries_0_rs2Val; // @[LSUQueue.scala 43:22]
  reg [7:0] entries_0_id; // @[LSUQueue.scala 43:22]
  reg [4:0] entries_0_rd; // @[LSUQueue.scala 43:22]
  reg  entries_1_busy; // @[LSUQueue.scala 43:22]
  reg  entries_1_ready; // @[LSUQueue.scala 43:22]
  reg  entries_1_decInfo_en; // @[LSUQueue.scala 43:22]
  reg  entries_1_decInfo_wen; // @[LSUQueue.scala 43:22]
  reg  entries_1_decInfo_load; // @[LSUQueue.scala 43:22]
  reg [1:0] entries_1_decInfo_wd; // @[LSUQueue.scala 43:22]
  reg  entries_1_decInfo_signed; // @[LSUQueue.scala 43:22]
  reg [31:0] entries_1_addr; // @[LSUQueue.scala 43:22]
  reg [31:0] entries_1_rs2Val; // @[LSUQueue.scala 43:22]
  reg [7:0] entries_1_id; // @[LSUQueue.scala 43:22]
  reg [4:0] entries_1_rd; // @[LSUQueue.scala 43:22]
  reg  entries_2_busy; // @[LSUQueue.scala 43:22]
  reg  entries_2_ready; // @[LSUQueue.scala 43:22]
  reg  entries_2_decInfo_en; // @[LSUQueue.scala 43:22]
  reg  entries_2_decInfo_wen; // @[LSUQueue.scala 43:22]
  reg  entries_2_decInfo_load; // @[LSUQueue.scala 43:22]
  reg [1:0] entries_2_decInfo_wd; // @[LSUQueue.scala 43:22]
  reg  entries_2_decInfo_signed; // @[LSUQueue.scala 43:22]
  reg [31:0] entries_2_addr; // @[LSUQueue.scala 43:22]
  reg [31:0] entries_2_rs2Val; // @[LSUQueue.scala 43:22]
  reg [7:0] entries_2_id; // @[LSUQueue.scala 43:22]
  reg [4:0] entries_2_rd; // @[LSUQueue.scala 43:22]
  reg  entries_3_busy; // @[LSUQueue.scala 43:22]
  reg  entries_3_ready; // @[LSUQueue.scala 43:22]
  reg  entries_3_decInfo_en; // @[LSUQueue.scala 43:22]
  reg  entries_3_decInfo_wen; // @[LSUQueue.scala 43:22]
  reg  entries_3_decInfo_load; // @[LSUQueue.scala 43:22]
  reg [1:0] entries_3_decInfo_wd; // @[LSUQueue.scala 43:22]
  reg  entries_3_decInfo_signed; // @[LSUQueue.scala 43:22]
  reg [31:0] entries_3_addr; // @[LSUQueue.scala 43:22]
  reg [31:0] entries_3_rs2Val; // @[LSUQueue.scala 43:22]
  reg [7:0] entries_3_id; // @[LSUQueue.scala 43:22]
  reg [4:0] entries_3_rd; // @[LSUQueue.scala 43:22]
  reg [1:0] head; // @[LSUQueue.scala 44:23]
  reg [1:0] tail; // @[LSUQueue.scala 45:23]
  reg [2:0] count; // @[LSUQueue.scala 47:24]
  wire  full = count == 3'h4; // @[LSUQueue.scala 48:22]
  wire  _GEN_1 = 2'h1 == tail ? entries_1_busy : entries_0_busy; // @[LSUQueue.scala 51:{30,30}]
  wire  _GEN_2 = 2'h2 == tail ? entries_2_busy : _GEN_1; // @[LSUQueue.scala 51:{30,30}]
  wire  _GEN_3 = 2'h3 == tail ? entries_3_busy : _GEN_2; // @[LSUQueue.scala 51:{30,30}]
  wire  _GEN_5 = 2'h1 == head ? entries_1_busy : entries_0_busy; // @[LSUQueue.scala 52:{40,40}]
  wire  _GEN_6 = 2'h2 == head ? entries_2_busy : _GEN_5; // @[LSUQueue.scala 52:{40,40}]
  wire  _GEN_7 = 2'h3 == head ? entries_3_busy : _GEN_6; // @[LSUQueue.scala 52:{40,40}]
  wire  _GEN_9 = 2'h1 == head ? entries_1_ready : entries_0_ready; // @[LSUQueue.scala 52:{40,40}]
  wire  _GEN_10 = 2'h2 == head ? entries_2_ready : _GEN_9; // @[LSUQueue.scala 52:{40,40}]
  wire  _GEN_11 = 2'h3 == head ? entries_3_ready : _GEN_10; // @[LSUQueue.scala 52:{40,40}]
  wire [31:0] _GEN_13 = 2'h1 == head ? entries_1_addr : entries_0_addr; // @[LSUQueue.scala 53:{22,22}]
  wire [31:0] _GEN_14 = 2'h2 == head ? entries_2_addr : _GEN_13; // @[LSUQueue.scala 53:{22,22}]
  wire  _GEN_17 = 2'h1 == head ? entries_1_decInfo_en : entries_0_decInfo_en; // @[LSUQueue.scala 54:{25,25}]
  wire  _GEN_18 = 2'h2 == head ? entries_2_decInfo_en : _GEN_17; // @[LSUQueue.scala 54:{25,25}]
  wire  _GEN_21 = 2'h1 == head ? entries_1_decInfo_wen : entries_0_decInfo_wen; // @[LSUQueue.scala 54:{25,25}]
  wire  _GEN_22 = 2'h2 == head ? entries_2_decInfo_wen : _GEN_21; // @[LSUQueue.scala 54:{25,25}]
  wire  _GEN_25 = 2'h1 == head ? entries_1_decInfo_load : entries_0_decInfo_load; // @[LSUQueue.scala 54:{25,25}]
  wire  _GEN_26 = 2'h2 == head ? entries_2_decInfo_load : _GEN_25; // @[LSUQueue.scala 54:{25,25}]
  wire [1:0] _GEN_29 = 2'h1 == head ? entries_1_decInfo_wd : entries_0_decInfo_wd; // @[LSUQueue.scala 54:{25,25}]
  wire [1:0] _GEN_30 = 2'h2 == head ? entries_2_decInfo_wd : _GEN_29; // @[LSUQueue.scala 54:{25,25}]
  wire  _GEN_33 = 2'h1 == head ? entries_1_decInfo_signed : entries_0_decInfo_signed; // @[LSUQueue.scala 54:{25,25}]
  wire  _GEN_34 = 2'h2 == head ? entries_2_decInfo_signed : _GEN_33; // @[LSUQueue.scala 54:{25,25}]
  wire [7:0] _GEN_37 = 2'h1 == head ? entries_1_id : entries_0_id; // @[LSUQueue.scala 55:{20,20}]
  wire [7:0] _GEN_38 = 2'h2 == head ? entries_2_id : _GEN_37; // @[LSUQueue.scala 55:{20,20}]
  wire [4:0] _GEN_41 = 2'h1 == head ? entries_1_rd : entries_0_rd; // @[LSUQueue.scala 56:{20,20}]
  wire [4:0] _GEN_42 = 2'h2 == head ? entries_2_rd : _GEN_41; // @[LSUQueue.scala 56:{20,20}]
  wire [31:0] _GEN_45 = 2'h1 == head ? entries_1_rs2Val : entries_0_rs2Val; // @[LSUQueue.scala 57:{24,24}]
  wire [31:0] _GEN_46 = 2'h2 == head ? entries_2_rs2Val : _GEN_45; // @[LSUQueue.scala 57:{24,24}]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_48 = 2'h0 == tail | entries_0_busy; // @[LSUQueue.scala 43:22 61:{28,28}]
  wire  _GEN_49 = 2'h1 == tail | entries_1_busy; // @[LSUQueue.scala 43:22 61:{28,28}]
  wire  _GEN_50 = 2'h2 == tail | entries_2_busy; // @[LSUQueue.scala 43:22 61:{28,28}]
  wire  _GEN_51 = 2'h3 == tail | entries_3_busy; // @[LSUQueue.scala 43:22 61:{28,28}]
  wire  _entries_ready_T = io_enq_bits_decInfo_wen ? 1'h0 : 1'h1; // @[LSUQueue.scala 67:35]
  wire  _GEN_88 = 2'h0 == tail ? _entries_ready_T : entries_0_ready; // @[LSUQueue.scala 43:22 67:{29,29}]
  wire  _GEN_89 = 2'h1 == tail ? _entries_ready_T : entries_1_ready; // @[LSUQueue.scala 43:22 67:{29,29}]
  wire  _GEN_90 = 2'h2 == tail ? _entries_ready_T : entries_2_ready; // @[LSUQueue.scala 43:22 67:{29,29}]
  wire  _GEN_91 = 2'h3 == tail ? _entries_ready_T : entries_3_ready; // @[LSUQueue.scala 43:22 67:{29,29}]
  wire [1:0] _tail_T_2 = tail + 2'h1; // @[LSUQueue.scala 69:60]
  wire  _GEN_92 = _T ? _GEN_48 : entries_0_busy; // @[LSUQueue.scala 43:22 59:24]
  wire  _GEN_93 = _T ? _GEN_49 : entries_1_busy; // @[LSUQueue.scala 43:22 59:24]
  wire  _GEN_94 = _T ? _GEN_50 : entries_2_busy; // @[LSUQueue.scala 43:22 59:24]
  wire  _GEN_95 = _T ? _GEN_51 : entries_3_busy; // @[LSUQueue.scala 43:22 59:24]
  wire  _GEN_132 = _T ? _GEN_88 : entries_0_ready; // @[LSUQueue.scala 43:22 59:24]
  wire  _GEN_133 = _T ? _GEN_89 : entries_1_ready; // @[LSUQueue.scala 43:22 59:24]
  wire  _GEN_134 = _T ? _GEN_90 : entries_2_ready; // @[LSUQueue.scala 43:22 59:24]
  wire  _GEN_135 = _T ? _GEN_91 : entries_3_ready; // @[LSUQueue.scala 43:22 59:24]
  wire  _T_1 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_141 = 2'h0 == head ? 1'h0 : _GEN_132; // @[LSUQueue.scala 74:{29,29}]
  wire  _GEN_142 = 2'h1 == head ? 1'h0 : _GEN_133; // @[LSUQueue.scala 74:{29,29}]
  wire  _GEN_143 = 2'h2 == head ? 1'h0 : _GEN_134; // @[LSUQueue.scala 74:{29,29}]
  wire  _GEN_144 = 2'h3 == head ? 1'h0 : _GEN_135; // @[LSUQueue.scala 74:{29,29}]
  wire [1:0] _head_T_2 = head + 2'h1; // @[LSUQueue.scala 76:60]
  wire  _GEN_149 = _T_1 ? _GEN_141 : _GEN_132; // @[LSUQueue.scala 72:24]
  wire  _GEN_150 = _T_1 ? _GEN_142 : _GEN_133; // @[LSUQueue.scala 72:24]
  wire  _GEN_151 = _T_1 ? _GEN_143 : _GEN_134; // @[LSUQueue.scala 72:24]
  wire  _GEN_152 = _T_1 ? _GEN_144 : _GEN_135; // @[LSUQueue.scala 72:24]
  wire [2:0] _count_T_1 = count + 3'h1; // @[LSUQueue.scala 81:28]
  wire [2:0] _GEN_154 = _T ? _count_T_1 : count; // @[LSUQueue.scala 80:27 81:19 47:24]
  wire [2:0] _count_T_3 = count - 3'h1; // @[LSUQueue.scala 84:28]
  wire  _GEN_157 = io_rob_bits_id == entries_0_id | _GEN_149; // @[LSUQueue.scala 92:62 93:29]
  wire  _GEN_160 = io_rob_bits_id == entries_1_id | _GEN_150; // @[LSUQueue.scala 92:62 93:29]
  wire  _GEN_163 = io_rob_bits_id == entries_2_id | _GEN_151; // @[LSUQueue.scala 92:62 93:29]
  wire  _GEN_166 = io_rob_bits_id == entries_3_id | _GEN_152; // @[LSUQueue.scala 92:62 93:29]
  assign io_enq_ready = ~full & ~_GEN_3; // @[LSUQueue.scala 51:27]
  assign io_deq_valid = _GEN_7 & _GEN_11; // @[LSUQueue.scala 52:40]
  assign io_deq_bits_decInfo_en = 2'h3 == head ? entries_3_decInfo_en : _GEN_18; // @[LSUQueue.scala 54:{25,25}]
  assign io_deq_bits_decInfo_wen = 2'h3 == head ? entries_3_decInfo_wen : _GEN_22; // @[LSUQueue.scala 54:{25,25}]
  assign io_deq_bits_decInfo_load = 2'h3 == head ? entries_3_decInfo_load : _GEN_26; // @[LSUQueue.scala 54:{25,25}]
  assign io_deq_bits_decInfo_wd = 2'h3 == head ? entries_3_decInfo_wd : _GEN_30; // @[LSUQueue.scala 54:{25,25}]
  assign io_deq_bits_decInfo_signed = 2'h3 == head ? entries_3_decInfo_signed : _GEN_34; // @[LSUQueue.scala 54:{25,25}]
  assign io_deq_bits_addr = 2'h3 == head ? entries_3_addr : _GEN_14; // @[LSUQueue.scala 53:{22,22}]
  assign io_deq_bits_rs2Val = 2'h3 == head ? entries_3_rs2Val : _GEN_46; // @[LSUQueue.scala 57:{24,24}]
  assign io_deq_bits_id = 2'h3 == head ? entries_3_id : _GEN_38; // @[LSUQueue.scala 55:{20,20}]
  assign io_deq_bits_rd = 2'h3 == head ? entries_3_rd : _GEN_42; // @[LSUQueue.scala 56:{20,20}]
  always @(posedge clock) begin
    if (io_flush) begin // @[LSUQueue.scala 99:21]
      entries_0_busy <= 1'h0; // @[LSUQueue.scala 100:37]
    end else if (_T_1) begin // @[LSUQueue.scala 72:24]
      if (2'h0 == head) begin // @[LSUQueue.scala 73:28]
        entries_0_busy <= 1'h0; // @[LSUQueue.scala 73:28]
      end else begin
        entries_0_busy <= _GEN_92;
      end
    end else begin
      entries_0_busy <= _GEN_92;
    end
    if (entries_0_busy) begin // @[LSUQueue.scala 89:22]
      if (~entries_0_ready) begin // @[LSUQueue.scala 90:28]
        entries_0_ready <= _GEN_157;
      end else begin
        entries_0_ready <= _GEN_149;
      end
    end else begin
      entries_0_ready <= _GEN_149;
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h0 == tail) begin // @[LSUQueue.scala 63:31]
        entries_0_decInfo_en <= io_enq_bits_decInfo_en; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h0 == tail) begin // @[LSUQueue.scala 63:31]
        entries_0_decInfo_wen <= io_enq_bits_decInfo_wen; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h0 == tail) begin // @[LSUQueue.scala 63:31]
        entries_0_decInfo_load <= io_enq_bits_decInfo_load; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h0 == tail) begin // @[LSUQueue.scala 63:31]
        entries_0_decInfo_wd <= io_enq_bits_decInfo_wd; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h0 == tail) begin // @[LSUQueue.scala 63:31]
        entries_0_decInfo_signed <= io_enq_bits_decInfo_signed; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h0 == tail) begin // @[LSUQueue.scala 62:28]
        entries_0_addr <= io_enq_bits_addr; // @[LSUQueue.scala 62:28]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h0 == tail) begin // @[LSUQueue.scala 66:30]
        entries_0_rs2Val <= io_enq_bits_rs2Val; // @[LSUQueue.scala 66:30]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h0 == tail) begin // @[LSUQueue.scala 64:26]
        entries_0_id <= io_enq_bits_id; // @[LSUQueue.scala 64:26]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h0 == tail) begin // @[LSUQueue.scala 65:26]
        entries_0_rd <= io_enq_bits_rd; // @[LSUQueue.scala 65:26]
      end
    end
    if (io_flush) begin // @[LSUQueue.scala 99:21]
      entries_1_busy <= 1'h0; // @[LSUQueue.scala 100:37]
    end else if (_T_1) begin // @[LSUQueue.scala 72:24]
      if (2'h1 == head) begin // @[LSUQueue.scala 73:28]
        entries_1_busy <= 1'h0; // @[LSUQueue.scala 73:28]
      end else begin
        entries_1_busy <= _GEN_93;
      end
    end else begin
      entries_1_busy <= _GEN_93;
    end
    if (entries_1_busy) begin // @[LSUQueue.scala 89:22]
      if (~entries_1_ready) begin // @[LSUQueue.scala 90:28]
        entries_1_ready <= _GEN_160;
      end else begin
        entries_1_ready <= _GEN_150;
      end
    end else begin
      entries_1_ready <= _GEN_150;
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h1 == tail) begin // @[LSUQueue.scala 63:31]
        entries_1_decInfo_en <= io_enq_bits_decInfo_en; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h1 == tail) begin // @[LSUQueue.scala 63:31]
        entries_1_decInfo_wen <= io_enq_bits_decInfo_wen; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h1 == tail) begin // @[LSUQueue.scala 63:31]
        entries_1_decInfo_load <= io_enq_bits_decInfo_load; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h1 == tail) begin // @[LSUQueue.scala 63:31]
        entries_1_decInfo_wd <= io_enq_bits_decInfo_wd; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h1 == tail) begin // @[LSUQueue.scala 63:31]
        entries_1_decInfo_signed <= io_enq_bits_decInfo_signed; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h1 == tail) begin // @[LSUQueue.scala 62:28]
        entries_1_addr <= io_enq_bits_addr; // @[LSUQueue.scala 62:28]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h1 == tail) begin // @[LSUQueue.scala 66:30]
        entries_1_rs2Val <= io_enq_bits_rs2Val; // @[LSUQueue.scala 66:30]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h1 == tail) begin // @[LSUQueue.scala 64:26]
        entries_1_id <= io_enq_bits_id; // @[LSUQueue.scala 64:26]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h1 == tail) begin // @[LSUQueue.scala 65:26]
        entries_1_rd <= io_enq_bits_rd; // @[LSUQueue.scala 65:26]
      end
    end
    if (io_flush) begin // @[LSUQueue.scala 99:21]
      entries_2_busy <= 1'h0; // @[LSUQueue.scala 100:37]
    end else if (_T_1) begin // @[LSUQueue.scala 72:24]
      if (2'h2 == head) begin // @[LSUQueue.scala 73:28]
        entries_2_busy <= 1'h0; // @[LSUQueue.scala 73:28]
      end else begin
        entries_2_busy <= _GEN_94;
      end
    end else begin
      entries_2_busy <= _GEN_94;
    end
    if (entries_2_busy) begin // @[LSUQueue.scala 89:22]
      if (~entries_2_ready) begin // @[LSUQueue.scala 90:28]
        entries_2_ready <= _GEN_163;
      end else begin
        entries_2_ready <= _GEN_151;
      end
    end else begin
      entries_2_ready <= _GEN_151;
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h2 == tail) begin // @[LSUQueue.scala 63:31]
        entries_2_decInfo_en <= io_enq_bits_decInfo_en; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h2 == tail) begin // @[LSUQueue.scala 63:31]
        entries_2_decInfo_wen <= io_enq_bits_decInfo_wen; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h2 == tail) begin // @[LSUQueue.scala 63:31]
        entries_2_decInfo_load <= io_enq_bits_decInfo_load; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h2 == tail) begin // @[LSUQueue.scala 63:31]
        entries_2_decInfo_wd <= io_enq_bits_decInfo_wd; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h2 == tail) begin // @[LSUQueue.scala 63:31]
        entries_2_decInfo_signed <= io_enq_bits_decInfo_signed; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h2 == tail) begin // @[LSUQueue.scala 62:28]
        entries_2_addr <= io_enq_bits_addr; // @[LSUQueue.scala 62:28]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h2 == tail) begin // @[LSUQueue.scala 66:30]
        entries_2_rs2Val <= io_enq_bits_rs2Val; // @[LSUQueue.scala 66:30]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h2 == tail) begin // @[LSUQueue.scala 64:26]
        entries_2_id <= io_enq_bits_id; // @[LSUQueue.scala 64:26]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h2 == tail) begin // @[LSUQueue.scala 65:26]
        entries_2_rd <= io_enq_bits_rd; // @[LSUQueue.scala 65:26]
      end
    end
    if (io_flush) begin // @[LSUQueue.scala 99:21]
      entries_3_busy <= 1'h0; // @[LSUQueue.scala 100:37]
    end else if (_T_1) begin // @[LSUQueue.scala 72:24]
      if (2'h3 == head) begin // @[LSUQueue.scala 73:28]
        entries_3_busy <= 1'h0; // @[LSUQueue.scala 73:28]
      end else begin
        entries_3_busy <= _GEN_95;
      end
    end else begin
      entries_3_busy <= _GEN_95;
    end
    if (entries_3_busy) begin // @[LSUQueue.scala 89:22]
      if (~entries_3_ready) begin // @[LSUQueue.scala 90:28]
        entries_3_ready <= _GEN_166;
      end else begin
        entries_3_ready <= _GEN_152;
      end
    end else begin
      entries_3_ready <= _GEN_152;
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h3 == tail) begin // @[LSUQueue.scala 63:31]
        entries_3_decInfo_en <= io_enq_bits_decInfo_en; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h3 == tail) begin // @[LSUQueue.scala 63:31]
        entries_3_decInfo_wen <= io_enq_bits_decInfo_wen; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h3 == tail) begin // @[LSUQueue.scala 63:31]
        entries_3_decInfo_load <= io_enq_bits_decInfo_load; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h3 == tail) begin // @[LSUQueue.scala 63:31]
        entries_3_decInfo_wd <= io_enq_bits_decInfo_wd; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h3 == tail) begin // @[LSUQueue.scala 63:31]
        entries_3_decInfo_signed <= io_enq_bits_decInfo_signed; // @[LSUQueue.scala 63:31]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h3 == tail) begin // @[LSUQueue.scala 62:28]
        entries_3_addr <= io_enq_bits_addr; // @[LSUQueue.scala 62:28]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h3 == tail) begin // @[LSUQueue.scala 66:30]
        entries_3_rs2Val <= io_enq_bits_rs2Val; // @[LSUQueue.scala 66:30]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h3 == tail) begin // @[LSUQueue.scala 64:26]
        entries_3_id <= io_enq_bits_id; // @[LSUQueue.scala 64:26]
      end
    end
    if (_T) begin // @[LSUQueue.scala 59:24]
      if (2'h3 == tail) begin // @[LSUQueue.scala 65:26]
        entries_3_rd <= io_enq_bits_rd; // @[LSUQueue.scala 65:26]
      end
    end
    if (reset) begin // @[LSUQueue.scala 44:23]
      head <= 2'h0; // @[LSUQueue.scala 44:23]
    end else if (io_flush) begin // @[LSUQueue.scala 99:21]
      head <= 2'h0; // @[LSUQueue.scala 101:14]
    end else if (_T_1) begin // @[LSUQueue.scala 72:24]
      if (head == 2'h3) begin // @[LSUQueue.scala 76:20]
        head <= 2'h0;
      end else begin
        head <= _head_T_2;
      end
    end
    if (reset) begin // @[LSUQueue.scala 45:23]
      tail <= 2'h0; // @[LSUQueue.scala 45:23]
    end else if (io_flush) begin // @[LSUQueue.scala 99:21]
      tail <= 2'h0; // @[LSUQueue.scala 102:14]
    end else if (_T) begin // @[LSUQueue.scala 59:24]
      if (tail == 2'h3) begin // @[LSUQueue.scala 69:20]
        tail <= 2'h0;
      end else begin
        tail <= _tail_T_2;
      end
    end
    if (reset) begin // @[LSUQueue.scala 47:24]
      count <= 3'h0; // @[LSUQueue.scala 47:24]
    end else if (io_flush) begin // @[LSUQueue.scala 99:21]
      count <= 3'h0; // @[LSUQueue.scala 103:15]
    end else if (~(_T_1 & _T)) begin // @[LSUQueue.scala 79:43]
      if (_T_1) begin // @[LSUQueue.scala 83:27]
        count <= _count_T_3; // @[LSUQueue.scala 84:19]
      end else begin
        count <= _GEN_154;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  entries_0_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  entries_0_ready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  entries_0_decInfo_en = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  entries_0_decInfo_wen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  entries_0_decInfo_load = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  entries_0_decInfo_wd = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  entries_0_decInfo_signed = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  entries_0_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  entries_0_rs2Val = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  entries_0_id = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  entries_0_rd = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  entries_1_busy = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  entries_1_ready = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  entries_1_decInfo_en = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  entries_1_decInfo_wen = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  entries_1_decInfo_load = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  entries_1_decInfo_wd = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  entries_1_decInfo_signed = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  entries_1_addr = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  entries_1_rs2Val = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  entries_1_id = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  entries_1_rd = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  entries_2_busy = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  entries_2_ready = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  entries_2_decInfo_en = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  entries_2_decInfo_wen = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  entries_2_decInfo_load = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  entries_2_decInfo_wd = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  entries_2_decInfo_signed = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  entries_2_addr = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  entries_2_rs2Val = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  entries_2_id = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  entries_2_rd = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  entries_3_busy = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  entries_3_ready = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  entries_3_decInfo_en = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  entries_3_decInfo_wen = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  entries_3_decInfo_load = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  entries_3_decInfo_wd = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  entries_3_decInfo_signed = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  entries_3_addr = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  entries_3_rs2Val = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  entries_3_id = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  entries_3_rd = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  head = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  tail = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  count = _RAND_46[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSUStage_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [4:0]  io_in_bits_lsuOp,
  input  [2:0]  io_in_bits_immSrc,
  input  [31:0] io_in_bits_rs1Val,
  input  [31:0] io_in_bits_rs2Val,
  input  [31:0] io_in_bits_inst,
  input  [7:0]  io_in_bits_id,
  output        io_out_valid,
  output [4:0]  io_out_bits_rd,
  output [31:0] io_out_bits_data,
  output [7:0]  io_out_bits_id,
  input         io_cache_read_req_ready,
  output        io_cache_read_req_valid,
  output [31:0] io_cache_read_req_bits_addr,
  output        io_cache_read_resp_ready,
  input         io_cache_read_resp_valid,
  input  [31:0] io_cache_read_resp_bits_data,
  input         io_cache_write_req_ready,
  output        io_cache_write_req_valid,
  output [31:0] io_cache_write_req_bits_addr,
  output [31:0] io_cache_write_req_bits_data,
  output [3:0]  io_cache_write_req_bits_mask,
  output        io_cache_write_resp_ready,
  input         io_cache_write_resp_valid,
  input  [7:0]  io_rob_bits_id,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  lsuQueue_clock; // @[LSU.scala 259:26]
  wire  lsuQueue_reset; // @[LSU.scala 259:26]
  wire  lsuQueue_io_enq_ready; // @[LSU.scala 259:26]
  wire  lsuQueue_io_enq_valid; // @[LSU.scala 259:26]
  wire  lsuQueue_io_enq_bits_decInfo_en; // @[LSU.scala 259:26]
  wire  lsuQueue_io_enq_bits_decInfo_wen; // @[LSU.scala 259:26]
  wire  lsuQueue_io_enq_bits_decInfo_load; // @[LSU.scala 259:26]
  wire [1:0] lsuQueue_io_enq_bits_decInfo_wd; // @[LSU.scala 259:26]
  wire  lsuQueue_io_enq_bits_decInfo_signed; // @[LSU.scala 259:26]
  wire [31:0] lsuQueue_io_enq_bits_addr; // @[LSU.scala 259:26]
  wire [31:0] lsuQueue_io_enq_bits_rs2Val; // @[LSU.scala 259:26]
  wire [7:0] lsuQueue_io_enq_bits_id; // @[LSU.scala 259:26]
  wire [4:0] lsuQueue_io_enq_bits_rd; // @[LSU.scala 259:26]
  wire  lsuQueue_io_deq_ready; // @[LSU.scala 259:26]
  wire  lsuQueue_io_deq_valid; // @[LSU.scala 259:26]
  wire  lsuQueue_io_deq_bits_decInfo_en; // @[LSU.scala 259:26]
  wire  lsuQueue_io_deq_bits_decInfo_wen; // @[LSU.scala 259:26]
  wire  lsuQueue_io_deq_bits_decInfo_load; // @[LSU.scala 259:26]
  wire [1:0] lsuQueue_io_deq_bits_decInfo_wd; // @[LSU.scala 259:26]
  wire  lsuQueue_io_deq_bits_decInfo_signed; // @[LSU.scala 259:26]
  wire [31:0] lsuQueue_io_deq_bits_addr; // @[LSU.scala 259:26]
  wire [31:0] lsuQueue_io_deq_bits_rs2Val; // @[LSU.scala 259:26]
  wire [7:0] lsuQueue_io_deq_bits_id; // @[LSU.scala 259:26]
  wire [4:0] lsuQueue_io_deq_bits_rd; // @[LSU.scala 259:26]
  wire [7:0] lsuQueue_io_rob_bits_id; // @[LSU.scala 259:26]
  wire  lsuQueue_io_flush; // @[LSU.scala 259:26]
  wire [31:0] immGen_io_inst; // @[LSU.scala 279:24]
  wire [2:0] immGen_io_immSrc; // @[LSU.scala 279:24]
  wire  immGen_io_immSign; // @[LSU.scala 279:24]
  wire [31:0] immGen_io_imm; // @[LSU.scala 279:24]
  reg  s0_full; // @[LSU.scala 268:26]
  reg [4:0] s0_info_lsuOp; // @[Reg.scala 19:16]
  wire  _s0_valid_T_1 = s0_info_lsuOp == 5'h14; // @[LSU.scala 295:75]
  wire  s0_valid = s0_full & (s0_info_lsuOp != 5'h14 | s0_info_lsuOp == 5'h14 & io_out_valid); // @[LSU.scala 295:25]
  wire  s0_fire = s0_valid & lsuQueue_io_enq_ready; // @[LSU.scala 269:28]
  wire  s0_ready = ~s0_full | s0_fire; // @[LSU.scala 274:26]
  wire  s0_latch = io_in_valid & s0_ready; // @[LSU.scala 267:32]
  reg [2:0] s0_info_immSrc; // @[Reg.scala 19:16]
  reg [31:0] s0_info_rs1Val; // @[Reg.scala 19:16]
  reg [31:0] s0_info_rs2Val; // @[Reg.scala 19:16]
  reg [31:0] s0_info_inst; // @[Reg.scala 19:16]
  reg [7:0] s0_info_id; // @[Reg.scala 19:16]
  wire [4:0] rd = s0_info_inst[11:7]; // @[util.scala 71:31]
  wire  _GEN_6 = s0_fire & s0_full ? 1'h0 : s0_full; // @[LSU.scala 268:26 277:{35,45}]
  wire  _GEN_7 = s0_latch | _GEN_6; // @[LSU.scala 276:{20,30}]
  wire  _T_2 = 5'h1 == s0_info_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_4 = 5'h2 == s0_info_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_6 = 5'h3 == s0_info_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_8 = 5'h4 == s0_info_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_10 = 5'h5 == s0_info_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_12 = 5'h6 == s0_info_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_14 = 5'h7 == s0_info_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_16 = 5'h8 == s0_info_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_31 = _T_10 ? 1'h0 : _T_12 | (_T_14 | _T_16); // @[Lookup.scala 34:39]
  wire  _T_32 = _T_8 ? 1'h0 : _T_31; // @[Lookup.scala 34:39]
  wire  _T_33 = _T_6 ? 1'h0 : _T_32; // @[Lookup.scala 34:39]
  wire  _T_34 = _T_4 ? 1'h0 : _T_33; // @[Lookup.scala 34:39]
  wire [1:0] _T_44 = _T_16 ? 2'h2 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _T_45 = _T_14 ? 2'h1 : _T_44; // @[Lookup.scala 34:39]
  wire [1:0] _T_46 = _T_12 ? 2'h0 : _T_45; // @[Lookup.scala 34:39]
  wire [1:0] _T_47 = _T_10 ? 2'h1 : _T_46; // @[Lookup.scala 34:39]
  wire [1:0] _T_48 = _T_8 ? 2'h0 : _T_47; // @[Lookup.scala 34:39]
  wire [1:0] _T_49 = _T_6 ? 2'h2 : _T_48; // @[Lookup.scala 34:39]
  wire [1:0] _T_50 = _T_4 ? 2'h1 : _T_49; // @[Lookup.scala 34:39]
  reg  s1_full; // @[LSU.scala 311:26]
  reg  s2_full; // @[LSU.scala 378:26]
  wire  _s2_loadRespValid_T = io_cache_read_resp_ready & io_cache_read_resp_valid; // @[Decoupled.scala 51:35]
  reg  s2_loadRespValid_holdReg; // @[Reg.scala 19:16]
  wire  s2_loadRespValid = _s2_loadRespValid_T ? io_cache_read_resp_valid : s2_loadRespValid_holdReg; // @[util.scala 26:12]
  wire  _s2_storeRespValid_T = io_cache_write_resp_ready & io_cache_write_resp_valid; // @[Decoupled.scala 51:35]
  reg  s2_storeRespValid_holdReg; // @[Reg.scala 19:16]
  wire  s2_storeRespValid = _s2_storeRespValid_T ? io_cache_write_resp_valid : s2_storeRespValid_holdReg; // @[util.scala 26:12]
  wire  s2_valid = s2_full & (s2_loadRespValid | s2_storeRespValid); // @[LSU.scala 413:25]
  wire  s2_fire = s2_valid & io_out_valid; // @[LSU.scala 379:28]
  wire  s2_ready = ~s2_full | s2_fire; // @[LSU.scala 387:26]
  wire  s1_ready = ~s1_full & s2_ready; // @[LSU.scala 320:30]
  wire  s1_latch = lsuQueue_io_deq_valid & s1_ready; // @[LSU.scala 310:42]
  wire  _s1_valid_T = io_cache_read_req_ready & io_cache_read_req_valid; // @[Decoupled.scala 51:35]
  wire  _s1_valid_T_1 = io_cache_write_req_ready & io_cache_write_req_valid; // @[Decoupled.scala 51:35]
  reg  s1_reqSend; // @[LSU.scala 347:29]
  wire  _s1_valid_T_3 = _s1_valid_T | _s1_valid_T_1 | s1_reqSend; // @[LSU.scala 371:79]
  wire  s1_valid = s1_full & (_s1_valid_T | _s1_valid_T_1 | s1_reqSend); // @[LSU.scala 371:25]
  wire  s1_fire = s1_valid & s2_ready; // @[LSU.scala 312:28]
  reg [4:0] s1_rd; // @[Reg.scala 19:16]
  reg [31:0] s1_rs2Val; // @[Reg.scala 19:16]
  reg [31:0] s1_addr; // @[Reg.scala 19:16]
  wire [1:0] s1_offset = s1_addr[1:0]; // @[LSU.scala 317:28]
  reg [7:0] s1_id; // @[Reg.scala 19:16]
  reg  s1_decInfo_en; // @[Reg.scala 19:16]
  reg  s1_decInfo_wen; // @[Reg.scala 19:16]
  reg  s1_decInfo_load; // @[Reg.scala 19:16]
  reg [1:0] s1_decInfo_wd; // @[Reg.scala 19:16]
  reg  s1_decInfo_signed; // @[Reg.scala 19:16]
  wire  _GEN_17 = s1_fire & s1_full ? 1'h0 : s1_full; // @[LSU.scala 311:26 324:{35,45}]
  wire  _GEN_18 = s1_latch | _GEN_17; // @[LSU.scala 323:{20,30}]
  wire  _io_cache_read_req_valid_T_1 = ~s1_reqSend; // @[LSU.scala 352:54]
  wire  _io_cache_read_req_valid_T_3 = ~io_flush; // @[LSU.scala 352:69]
  wire [4:0] _io_cache_write_req_bits_data_T = {s1_offset, 3'h0}; // @[LSU.scala 357:60]
  wire [62:0] _GEN_0 = {{31'd0}, s1_rs2Val}; // @[LSU.scala 357:46]
  wire [62:0] _io_cache_write_req_bits_data_T_1 = _GEN_0 << _io_cache_write_req_bits_data_T; // @[LSU.scala 357:46]
  wire [3:0] _s1_storeMask_T_1 = 4'h1 << s1_offset; // @[OneHot.scala 57:35]
  wire [2:0] _s1_storeMask_T_6 = 2'h1 == s1_offset ? 3'h6 : 3'h3; // @[Mux.scala 81:58]
  wire [3:0] _s1_storeMask_T_8 = 2'h2 == s1_offset ? 4'hc : {{1'd0}, _s1_storeMask_T_6}; // @[Mux.scala 81:58]
  wire [3:0] _s1_storeMask_T_10 = 2'h0 == s1_decInfo_wd ? _s1_storeMask_T_1 : 4'hf; // @[Mux.scala 81:58]
  wire [3:0] _s1_storeMask_T_12 = 2'h1 == s1_decInfo_wd ? _s1_storeMask_T_8 : _s1_storeMask_T_10; // @[Mux.scala 81:58]
  reg [4:0] s2_rd; // @[Reg.scala 19:16]
  reg  s2_load; // @[Reg.scala 19:16]
  reg  s2_en; // @[Reg.scala 19:16]
  reg  s2_signed; // @[Reg.scala 19:16]
  reg [1:0] s2_width; // @[Reg.scala 19:16]
  reg [1:0] s2_offset; // @[Reg.scala 19:16]
  reg [7:0] s2_id; // @[Reg.scala 19:16]
  wire  _GEN_28 = s2_fire & s2_full ? 1'h0 : s2_full; // @[LSU.scala 378:26 390:{35,45}]
  wire  _GEN_29 = s1_fire | _GEN_28; // @[LSU.scala 389:{20,30}]
  reg [31:0] s2_loadResp_holdReg_data; // @[Reg.scala 19:16]
  wire [31:0] _GEN_30 = _s2_loadRespValid_T ? io_cache_read_resp_bits_data : s2_loadResp_holdReg_data; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _s2_loadDataRaw_T_2 = {8'h0,_GEN_30[31:8]}; // @[Cat.scala 33:92]
  wire [31:0] _s2_loadDataRaw_T_5 = {16'h0,_GEN_30[31:16]}; // @[Cat.scala 33:92]
  wire [31:0] _s2_loadDataRaw_T_8 = {24'h0,_GEN_30[31:24]}; // @[Cat.scala 33:92]
  wire [31:0] _s2_loadDataRaw_T_10 = 2'h1 == s2_offset ? _s2_loadDataRaw_T_2 : _GEN_30; // @[Mux.scala 81:58]
  wire [31:0] _s2_loadDataRaw_T_12 = 2'h2 == s2_offset ? _s2_loadDataRaw_T_5 : _s2_loadDataRaw_T_10; // @[Mux.scala 81:58]
  wire [31:0] s2_loadDataRaw = 2'h3 == s2_offset ? _s2_loadDataRaw_T_8 : _s2_loadDataRaw_T_12; // @[Mux.scala 81:58]
  wire [7:0] _s2_loadData_T_1 = s2_loadDataRaw[7:0]; // @[LSU.scala 407:88]
  wire  s2_loadData_signBit = _s2_loadData_T_1[7]; // @[util.scala 42:27]
  wire [5:0] s2_loadData_out_lo_lo = {s2_loadData_signBit,s2_loadData_signBit,s2_loadData_signBit,s2_loadData_signBit,
    s2_loadData_signBit,s2_loadData_signBit}; // @[Cat.scala 33:92]
  wire [11:0] s2_loadData_out_lo = {s2_loadData_signBit,s2_loadData_signBit,s2_loadData_signBit,s2_loadData_signBit,
    s2_loadData_signBit,s2_loadData_signBit,s2_loadData_out_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] _s2_loadData_out_T_1 = s2_loadDataRaw[7:0]; // @[util.scala 46:75]
  wire [31:0] s2_loadData_out = {s2_loadData_signBit,s2_loadData_signBit,s2_loadData_signBit,s2_loadData_signBit,
    s2_loadData_signBit,s2_loadData_signBit,s2_loadData_out_lo_lo,s2_loadData_out_lo,_s2_loadData_out_T_1}; // @[Cat.scala 33:92]
  wire [31:0] s2_loadData_out_1 = {{24'd0}, s2_loadDataRaw[7:0]}; // @[util.scala 62:36]
  wire [31:0] _s2_loadData_T_3 = s2_signed ? s2_loadData_out : s2_loadData_out_1; // @[LSU.scala 407:48]
  wire [15:0] _s2_loadData_T_5 = s2_loadDataRaw[15:0]; // @[LSU.scala 408:89]
  wire  s2_loadData_signBit_1 = _s2_loadData_T_5[15]; // @[util.scala 42:27]
  wire [7:0] s2_loadData_out_lo_1 = {s2_loadData_signBit_1,s2_loadData_signBit_1,s2_loadData_signBit_1,
    s2_loadData_signBit_1,s2_loadData_signBit_1,s2_loadData_signBit_1,s2_loadData_signBit_1,s2_loadData_signBit_1}; // @[Cat.scala 33:92]
  wire [15:0] _s2_loadData_out_T_3 = s2_loadDataRaw[15:0]; // @[util.scala 46:75]
  wire [31:0] s2_loadData_out_2 = {s2_loadData_signBit_1,s2_loadData_signBit_1,s2_loadData_signBit_1,
    s2_loadData_signBit_1,s2_loadData_signBit_1,s2_loadData_signBit_1,s2_loadData_signBit_1,s2_loadData_signBit_1,
    s2_loadData_out_lo_1,_s2_loadData_out_T_3}; // @[Cat.scala 33:92]
  wire [31:0] s2_loadData_out_3 = {{16'd0}, s2_loadDataRaw[15:0]}; // @[util.scala 62:36]
  wire [31:0] _s2_loadData_T_7 = s2_signed ? s2_loadData_out_2 : s2_loadData_out_3; // @[LSU.scala 408:48]
  wire [31:0] _s2_loadData_T_10 = 2'h3 == s2_offset ? _s2_loadDataRaw_T_8 : _s2_loadDataRaw_T_12; // @[util.scala 44:18]
  wire [31:0] _s2_loadData_T_12 = s2_signed ? _s2_loadData_T_10 : s2_loadDataRaw; // @[LSU.scala 409:48]
  wire [31:0] _s2_loadData_T_14 = 2'h0 == s2_width ? _s2_loadData_T_3 : s2_loadDataRaw; // @[Mux.scala 81:58]
  wire [31:0] _s2_loadData_T_16 = 2'h1 == s2_width ? _s2_loadData_T_7 : _s2_loadData_T_14; // @[Mux.scala 81:58]
  wire  s0_fence = s0_full & _s0_valid_T_1; // @[LSU.scala 415:28]
  LSUQueue lsuQueue ( // @[LSU.scala 259:26]
    .clock(lsuQueue_clock),
    .reset(lsuQueue_reset),
    .io_enq_ready(lsuQueue_io_enq_ready),
    .io_enq_valid(lsuQueue_io_enq_valid),
    .io_enq_bits_decInfo_en(lsuQueue_io_enq_bits_decInfo_en),
    .io_enq_bits_decInfo_wen(lsuQueue_io_enq_bits_decInfo_wen),
    .io_enq_bits_decInfo_load(lsuQueue_io_enq_bits_decInfo_load),
    .io_enq_bits_decInfo_wd(lsuQueue_io_enq_bits_decInfo_wd),
    .io_enq_bits_decInfo_signed(lsuQueue_io_enq_bits_decInfo_signed),
    .io_enq_bits_addr(lsuQueue_io_enq_bits_addr),
    .io_enq_bits_rs2Val(lsuQueue_io_enq_bits_rs2Val),
    .io_enq_bits_id(lsuQueue_io_enq_bits_id),
    .io_enq_bits_rd(lsuQueue_io_enq_bits_rd),
    .io_deq_ready(lsuQueue_io_deq_ready),
    .io_deq_valid(lsuQueue_io_deq_valid),
    .io_deq_bits_decInfo_en(lsuQueue_io_deq_bits_decInfo_en),
    .io_deq_bits_decInfo_wen(lsuQueue_io_deq_bits_decInfo_wen),
    .io_deq_bits_decInfo_load(lsuQueue_io_deq_bits_decInfo_load),
    .io_deq_bits_decInfo_wd(lsuQueue_io_deq_bits_decInfo_wd),
    .io_deq_bits_decInfo_signed(lsuQueue_io_deq_bits_decInfo_signed),
    .io_deq_bits_addr(lsuQueue_io_deq_bits_addr),
    .io_deq_bits_rs2Val(lsuQueue_io_deq_bits_rs2Val),
    .io_deq_bits_id(lsuQueue_io_deq_bits_id),
    .io_deq_bits_rd(lsuQueue_io_deq_bits_rd),
    .io_rob_bits_id(lsuQueue_io_rob_bits_id),
    .io_flush(lsuQueue_io_flush)
  );
  ImmGen immGen ( // @[LSU.scala 279:24]
    .io_inst(immGen_io_inst),
    .io_immSrc(immGen_io_immSrc),
    .io_immSign(immGen_io_immSign),
    .io_imm(immGen_io_imm)
  );
  assign io_in_ready = ~s0_full | s0_fire; // @[LSU.scala 274:26]
  assign io_out_valid = s2_valid & s2_en | s0_fence; // @[LSU.scala 416:39]
  assign io_out_bits_rd = s2_rd; // @[LSU.scala 417:20]
  assign io_out_bits_data = 2'h2 == s2_width ? _s2_loadData_T_12 : _s2_loadData_T_16; // @[Mux.scala 81:58]
  assign io_out_bits_id = s0_fence ? s0_info_id : s2_id; // @[LSU.scala 419:26]
  assign io_cache_read_req_valid = s1_decInfo_load & s1_full & ~s1_reqSend & ~io_flush; // @[LSU.scala 352:66]
  assign io_cache_read_req_bits_addr = {s1_addr[31:2],2'h0}; // @[Cat.scala 33:92]
  assign io_cache_read_resp_ready = s2_load; // @[LSU.scala 392:30]
  assign io_cache_write_req_valid = s1_decInfo_wen & s1_full & _io_cache_read_req_valid_T_1 &
    _io_cache_read_req_valid_T_3; // @[LSU.scala 355:66]
  assign io_cache_write_req_bits_addr = {s1_addr[31:2],2'h0}; // @[Cat.scala 33:92]
  assign io_cache_write_req_bits_data = _io_cache_write_req_bits_data_T_1[31:0]; // @[LSU.scala 357:34]
  assign io_cache_write_req_bits_mask = 2'h2 == s1_decInfo_wd ? 4'hf : _s1_storeMask_T_12; // @[Mux.scala 81:58]
  assign io_cache_write_resp_ready = ~s2_load; // @[LSU.scala 393:34]
  assign lsuQueue_clock = clock;
  assign lsuQueue_reset = reset;
  assign lsuQueue_io_enq_valid = s0_full & (s0_info_lsuOp != 5'h14 | s0_info_lsuOp == 5'h14 & io_out_valid); // @[LSU.scala 295:25]
  assign lsuQueue_io_enq_bits_decInfo_en = _T_2 | (_T_4 | (_T_6 | (_T_8 | (_T_10 | (_T_12 | (_T_14 | _T_16)))))); // @[Lookup.scala 34:39]
  assign lsuQueue_io_enq_bits_decInfo_wen = _T_2 ? 1'h0 : _T_34; // @[Lookup.scala 34:39]
  assign lsuQueue_io_enq_bits_decInfo_load = _T_2 | (_T_4 | (_T_6 | (_T_8 | _T_10))); // @[Lookup.scala 34:39]
  assign lsuQueue_io_enq_bits_decInfo_wd = _T_2 ? 2'h0 : _T_50; // @[Lookup.scala 34:39]
  assign lsuQueue_io_enq_bits_decInfo_signed = _T_2 | (_T_4 | (_T_6 | _T_32)); // @[Lookup.scala 34:39]
  assign lsuQueue_io_enq_bits_addr = immGen_io_imm + s0_info_rs1Val; // @[LSU.scala 281:26]
  assign lsuQueue_io_enq_bits_rs2Val = s0_info_rs2Val; // @[LSU.scala 303:33]
  assign lsuQueue_io_enq_bits_id = s0_info_id; // @[LSU.scala 301:29]
  assign lsuQueue_io_enq_bits_rd = s0_info_lsuOp == 5'h8 | s0_info_lsuOp == 5'h7 | s0_info_lsuOp == 5'h6 | _s0_valid_T_1
     ? 5'h0 : rd; // @[LSU.scala 273:20]
  assign lsuQueue_io_deq_ready = ~s1_full & s2_ready; // @[LSU.scala 320:30]
  assign lsuQueue_io_rob_bits_id = io_rob_bits_id; // @[LSU.scala 260:21]
  assign lsuQueue_io_flush = io_flush; // @[LSU.scala 261:23]
  assign immGen_io_inst = s0_info_inst; // @[LSU.scala 284:20]
  assign immGen_io_immSrc = s0_info_immSrc; // @[LSU.scala 282:22]
  assign immGen_io_immSign = 1'h1; // @[LSU.scala 283:23]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 268:26]
      s0_full <= 1'h0; // @[LSU.scala 268:26]
    end else if (io_flush) begin // @[LSU.scala 422:20]
      s0_full <= 1'h0; // @[LSU.scala 423:17]
    end else begin
      s0_full <= _GEN_7;
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_lsuOp <= io_in_bits_lsuOp; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_immSrc <= io_in_bits_immSrc; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_rs1Val <= io_in_bits_rs1Val; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_rs2Val <= io_in_bits_rs2Val; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_inst <= io_in_bits_inst; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_id <= io_in_bits_id; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[LSU.scala 311:26]
      s1_full <= 1'h0; // @[LSU.scala 311:26]
    end else if (io_flush) begin // @[LSU.scala 422:20]
      s1_full <= 1'h0; // @[LSU.scala 424:17]
    end else begin
      s1_full <= _GEN_18;
    end
    if (reset) begin // @[LSU.scala 378:26]
      s2_full <= 1'h0; // @[LSU.scala 378:26]
    end else if (io_flush) begin // @[LSU.scala 422:20]
      s2_full <= 1'h0; // @[LSU.scala 425:17]
    end else begin
      s2_full <= _GEN_29;
    end
    if (s1_fire) begin // @[util.scala 25:21]
      s2_loadRespValid_holdReg <= 1'h0; // @[util.scala 25:31]
    end else if (_s2_loadRespValid_T) begin // @[util.scala 26:12]
      s2_loadRespValid_holdReg <= io_cache_read_resp_valid;
    end
    if (s1_fire) begin // @[util.scala 25:21]
      s2_storeRespValid_holdReg <= 1'h0; // @[util.scala 25:31]
    end else if (_s2_storeRespValid_T) begin // @[util.scala 26:12]
      s2_storeRespValid_holdReg <= io_cache_write_resp_valid;
    end
    if (reset) begin // @[LSU.scala 347:29]
      s1_reqSend <= 1'h0; // @[LSU.scala 347:29]
    end else if (s1_fire) begin // @[LSU.scala 348:19]
      s1_reqSend <= 1'h0; // @[LSU.scala 348:32]
    end else begin
      s1_reqSend <= _s1_valid_T_3;
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_rd <= lsuQueue_io_deq_bits_rd; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_rs2Val <= lsuQueue_io_deq_bits_rs2Val; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_addr <= lsuQueue_io_deq_bits_addr; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_id <= lsuQueue_io_deq_bits_id; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_decInfo_en <= lsuQueue_io_deq_bits_decInfo_en; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_decInfo_wen <= lsuQueue_io_deq_bits_decInfo_wen; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_decInfo_load <= lsuQueue_io_deq_bits_decInfo_load; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_decInfo_wd <= lsuQueue_io_deq_bits_decInfo_wd; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_decInfo_signed <= lsuQueue_io_deq_bits_decInfo_signed; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_rd <= s1_rd; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_load <= s1_decInfo_load; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_en <= s1_decInfo_en; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_signed <= s1_decInfo_signed; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_width <= s1_decInfo_wd; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_offset <= s1_offset; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_id <= s1_id; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[util.scala 25:21]
      s2_loadResp_holdReg_data <= 32'h0; // @[util.scala 25:31]
    end else if (_s2_loadRespValid_T) begin // @[Reg.scala 20:18]
      s2_loadResp_holdReg_data <= io_cache_read_resp_bits_data; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s0_info_lsuOp = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  s0_info_immSrc = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  s0_info_rs1Val = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  s0_info_rs2Val = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  s0_info_inst = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  s0_info_id = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  s1_full = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s2_full = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  s2_loadRespValid_holdReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  s2_storeRespValid_holdReg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  s1_reqSend = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  s1_rd = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  s1_rs2Val = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  s1_addr = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  s1_id = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  s1_decInfo_en = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  s1_decInfo_wen = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  s1_decInfo_load = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  s1_decInfo_wd = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  s1_decInfo_signed = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  s2_rd = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  s2_load = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  s2_en = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  s2_signed = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  s2_width = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  s2_offset = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  s2_id = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  s2_loadResp_holdReg_data = _RAND_28[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CsrFile(
  input         clock,
  input         reset,
  input  [2:0]  io_read_op,
  output        io_read_valid,
  input  [11:0] io_read_addr,
  output [31:0] io_read_data,
  input  [2:0]  io_write_op,
  input  [11:0] io_write_addr,
  input  [31:0] io_write_data,
  output [31:0] io_mepc,
  output [31:0] io_trapVec,
  output [31:0] csrState_0_mcycle,
  output [31:0] csrState_0_mcycleh
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg  mcause_int; // @[CsrFile.scala 69:28]
  reg [30:0] mcause_code; // @[CsrFile.scala 69:28]
  reg  mstatus_sum; // @[CsrFile.scala 70:28]
  reg [1:0] mstatus_mpp; // @[CsrFile.scala 70:28]
  reg  mstatus_spp; // @[CsrFile.scala 70:28]
  reg  mstatus_mpie; // @[CsrFile.scala 70:28]
  reg  mstatus_spie; // @[CsrFile.scala 70:28]
  reg  mstatus_mie; // @[CsrFile.scala 70:28]
  reg  mstatus_sie; // @[CsrFile.scala 70:28]
  reg [29:0] mtvec_base; // @[CsrFile.scala 71:28]
  reg [1:0] mtvec_mode; // @[CsrFile.scala 71:28]
  reg [31:0] medeleg_data; // @[CsrFile.scala 72:28]
  reg [31:0] mideleg_data; // @[CsrFile.scala 73:28]
  reg [31:0] mepc_data; // @[CsrFile.scala 74:28]
  reg  satp_mode; // @[CsrFile.scala 75:28]
  reg [21:0] satp_ppn; // @[CsrFile.scala 75:28]
  reg [63:0] mcycle_data; // @[CsrFile.scala 77:28]
  wire [31:0] _T = {mcause_int,mcause_code}; // @[CsrFile.scala 88:49]
  wire [10:0] lo = {2'h0,mstatus_spp,mstatus_mpie,1'h0,mstatus_spie,1'h0,mstatus_mie,1'h0,mstatus_sie,1'h0}; // @[CsrFile.scala 89:50]
  wire [31:0] _T_1 = {13'h0,mstatus_sum,1'h0,2'h0,2'h0,mstatus_mpp,lo}; // @[CsrFile.scala 89:50]
  wire [31:0] _T_2 = {mtvec_base,mtvec_mode}; // @[CsrFile.scala 90:48]
  wire [31:0] _T_3 = {satp_mode,9'h0,satp_ppn}; // @[CsrFile.scala 94:47]
  wire  _T_7 = 12'hf14 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_9 = 12'h342 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_13 = 12'h305 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_15 = 12'h302 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_17 = 12'h303 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_19 = 12'h341 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_21 = 12'h180 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_23 = 12'h343 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_25 = 12'hb00 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_27 = 12'hb80 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_29 = 12'h3a0 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_31 = 12'h3a1 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_33 = 12'h3a2 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_35 = 12'h3a3 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_37 = 12'h3b0 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_39 = 12'h3b1 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_41 = 12'h3b2 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_43 = 12'h3b3 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_45 = 12'h3b4 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_47 = 12'h3b5 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_49 = 12'h3b6 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_51 = 12'h3b7 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_53 = 12'h3b8 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_55 = 12'h3b9 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_57 = 12'h3ba == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_59 = 12'h3bb == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_61 = 12'h3bc == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_63 = 12'h3bd == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_65 = 12'h3be == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_67 = 12'h3bf == io_read_addr; // @[Lookup.scala 31:38]
  wire [31:0] _T_88 = _T_27 ? mcycle_data[63:32] : 32'h0; // @[Lookup.scala 34:39]
  wire [31:0] _T_89 = _T_25 ? mcycle_data[31:0] : _T_88; // @[Lookup.scala 34:39]
  wire [31:0] _T_90 = _T_23 ? 32'h0 : _T_89; // @[Lookup.scala 34:39]
  wire [31:0] _T_91 = _T_21 ? _T_3 : _T_90; // @[Lookup.scala 34:39]
  wire [31:0] _T_92 = _T_19 ? mepc_data : _T_91; // @[Lookup.scala 34:39]
  wire [31:0] _T_93 = _T_17 ? mideleg_data : _T_92; // @[Lookup.scala 34:39]
  wire [31:0] _T_94 = _T_15 ? medeleg_data : _T_93; // @[Lookup.scala 34:39]
  wire [31:0] _T_95 = _T_13 ? _T_2 : _T_94; // @[Lookup.scala 34:39]
  wire [31:0] _T_96 = _T_9 ? _T_1 : _T_95; // @[Lookup.scala 34:39]
  wire [31:0] _T_97 = _T_9 ? _T : _T_96; // @[Lookup.scala 34:39]
  wire  readable = _T_7 | (_T_9 | (_T_9 | (_T_13 | (_T_15 | (_T_17 | (_T_19 | (_T_21 | (_T_23 | (_T_25 | (_T_27 | (_T_29
     | (_T_31 | (_T_33 | (_T_35 | (_T_37 | (_T_39 | (_T_41 | (_T_43 | (_T_45 | (_T_47 | (_T_49 | (_T_51 | (_T_53 | (
    _T_55 | (_T_57 | (_T_59 | (_T_61 | (_T_63 | (_T_65 | _T_67))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  writable = _T_7 ? 1'h0 : _T_9 | (_T_9 | (_T_13 | (_T_15 | (_T_17 | (_T_19 | (_T_21 | (_T_23 | (_T_25 | (_T_27 |
    (_T_29 | (_T_31 | (_T_33 | (_T_35 | (_T_37 | (_T_39 | (_T_41 | (_T_43 | (_T_45 | (_T_47 | (_T_49 | (_T_51 | (_T_53
     | (_T_55 | (_T_57 | (_T_59 | (_T_61 | (_T_63 | (_T_65 | _T_67)))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _readValid_T = readable & writable; // @[CsrFile.scala 130:30]
  wire  _readValid_T_6 = 3'h2 == io_read_op ? writable : 3'h1 == io_read_op & readable; // @[Mux.scala 81:58]
  wire  _readValid_T_8 = 3'h3 == io_read_op ? _readValid_T : _readValid_T_6; // @[Mux.scala 81:58]
  wire  _readValid_T_10 = 3'h4 == io_read_op ? _readValid_T : _readValid_T_8; // @[Mux.scala 81:58]
  wire  _csrData_T_1 = 12'hf14 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_3 = 12'h342 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_7 = 12'h305 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_9 = 12'h302 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_11 = 12'h303 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_13 = 12'h341 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_15 = 12'h180 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_17 = 12'h343 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_19 = 12'hb00 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_21 = 12'hb80 == io_write_addr; // @[Lookup.scala 31:38]
  wire [31:0] _csrData_T_82 = _csrData_T_21 ? mcycle_data[63:32] : 32'h0; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_83 = _csrData_T_19 ? mcycle_data[31:0] : _csrData_T_82; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_84 = _csrData_T_17 ? 32'h0 : _csrData_T_83; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_85 = _csrData_T_15 ? _T_3 : _csrData_T_84; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_86 = _csrData_T_13 ? mepc_data : _csrData_T_85; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_87 = _csrData_T_11 ? mideleg_data : _csrData_T_86; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_88 = _csrData_T_9 ? medeleg_data : _csrData_T_87; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_89 = _csrData_T_7 ? _T_2 : _csrData_T_88; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_90 = _csrData_T_3 ? _T_1 : _csrData_T_89; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_91 = _csrData_T_3 ? _T : _csrData_T_90; // @[Lookup.scala 34:39]
  wire [31:0] csrData = _csrData_T_1 ? 32'h0 : _csrData_T_91; // @[Lookup.scala 34:39]
  wire  writeEn = io_write_op != 3'h0 & io_write_op != 3'h1; // @[CsrFile.scala 140:43]
  wire [31:0] _writeData_T = csrData | io_write_data; // @[CsrFile.scala 144:29]
  wire [31:0] _writeData_T_1 = ~io_write_data; // @[CsrFile.scala 145:31]
  wire [31:0] _writeData_T_2 = csrData & _writeData_T_1; // @[CsrFile.scala 145:29]
  wire [31:0] _writeData_T_4 = 3'h2 == io_write_op ? io_write_data : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _writeData_T_6 = 3'h3 == io_write_op ? io_write_data : _writeData_T_4; // @[Mux.scala 81:58]
  wire [31:0] _writeData_T_8 = 3'h4 == io_write_op ? _writeData_T : _writeData_T_6; // @[Mux.scala 81:58]
  wire [31:0] writeData = 3'h5 == io_write_op ? _writeData_T_2 : _writeData_T_8; // @[Mux.scala 81:58]
  wire [63:0] _mcycle_data_T_1 = mcycle_data + 64'h1; // @[CsrFile.scala 148:32]
  wire [6:0] medeleg_data_lo = {writeData[6],1'h0,writeData[4:2],1'h0,writeData[0]}; // @[Cat.scala 33:92]
  wire [15:0] _medeleg_data_T_6 = {writeData[15],1'h0,writeData[13:12],2'h0,writeData[9:8],1'h0,medeleg_data_lo}; // @[Cat.scala 33:92]
  wire [11:0] _mideleg_data_T_3 = {2'h0,writeData[9],3'h0,writeData[5],3'h0,writeData[1],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] _mepc_data_T_1 = {writeData[31:2],2'h0}; // @[Cat.scala 33:92]
  wire [63:0] _mcycle_data_T_3 = {mcycle_data[63:32],writeData}; // @[Cat.scala 33:92]
  wire [63:0] _mcycle_data_T_5 = {writeData,mcycle_data[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_0 = _csrData_T_21 ? _mcycle_data_T_5 : _mcycle_data_T_1; // @[CsrFile.scala 148:17 151:31 160:43]
  wire [63:0] _GEN_1 = _csrData_T_19 ? _mcycle_data_T_3 : _GEN_0; // @[CsrFile.scala 151:31 159:43]
  wire  _GEN_2 = _csrData_T_15 ? writeData[31] : satp_mode; // @[CsrFile.scala 151:31 CSR.scala 187:11 CsrFile.scala 75:28]
  wire [21:0] _GEN_3 = _csrData_T_15 ? writeData[21:0] : satp_ppn; // @[CsrFile.scala 151:31 CSR.scala 188:11 CsrFile.scala 75:28]
  wire [63:0] _GEN_4 = _csrData_T_15 ? _mcycle_data_T_1 : _GEN_1; // @[CsrFile.scala 148:17 151:31]
  wire [31:0] _GEN_5 = _csrData_T_13 ? _mepc_data_T_1 : mepc_data; // @[CsrFile.scala 151:31 CSR.scala 369:11 CsrFile.scala 74:28]
  wire  _GEN_6 = _csrData_T_13 ? satp_mode : _GEN_2; // @[CsrFile.scala 151:31 75:28]
  wire [21:0] _GEN_7 = _csrData_T_13 ? satp_ppn : _GEN_3; // @[CsrFile.scala 151:31 75:28]
  wire [63:0] _GEN_8 = _csrData_T_13 ? _mcycle_data_T_1 : _GEN_4; // @[CsrFile.scala 148:17 151:31]
  wire [31:0] _GEN_9 = _csrData_T_11 ? {{20'd0}, _mideleg_data_T_3} : mideleg_data; // @[CsrFile.scala 151:31 CSR.scala 271:11 CsrFile.scala 73:28]
  wire [31:0] _GEN_10 = _csrData_T_11 ? mepc_data : _GEN_5; // @[CsrFile.scala 151:31 74:28]
  wire  _GEN_11 = _csrData_T_11 ? satp_mode : _GEN_6; // @[CsrFile.scala 151:31 75:28]
  wire [21:0] _GEN_12 = _csrData_T_11 ? satp_ppn : _GEN_7; // @[CsrFile.scala 151:31 75:28]
  wire [63:0] _GEN_13 = _csrData_T_11 ? _mcycle_data_T_1 : _GEN_8; // @[CsrFile.scala 148:17 151:31]
  wire [31:0] _GEN_14 = _csrData_T_9 ? {{16'd0}, _medeleg_data_T_6} : medeleg_data; // @[CsrFile.scala 151:31 CSR.scala 256:11 CsrFile.scala 72:28]
  wire [31:0] _GEN_15 = _csrData_T_9 ? mideleg_data : _GEN_9; // @[CsrFile.scala 151:31 73:28]
  wire [31:0] _GEN_16 = _csrData_T_9 ? mepc_data : _GEN_10; // @[CsrFile.scala 151:31 74:28]
  wire  _GEN_17 = _csrData_T_9 ? satp_mode : _GEN_11; // @[CsrFile.scala 151:31 75:28]
  wire [21:0] _GEN_18 = _csrData_T_9 ? satp_ppn : _GEN_12; // @[CsrFile.scala 151:31 75:28]
  wire [63:0] _GEN_19 = _csrData_T_9 ? _mcycle_data_T_1 : _GEN_13; // @[CsrFile.scala 148:17 151:31]
  wire [29:0] _GEN_20 = _csrData_T_7 ? writeData[31:2] : mtvec_base; // @[CsrFile.scala 151:31 CSR.scala 345:11 CsrFile.scala 71:28]
  wire [1:0] _GEN_21 = _csrData_T_7 ? {{1'd0}, writeData[0]} : mtvec_mode; // @[CsrFile.scala 151:31 CSR.scala 346:11 CsrFile.scala 71:28]
  wire [31:0] _GEN_22 = _csrData_T_7 ? medeleg_data : _GEN_14; // @[CsrFile.scala 151:31 72:28]
  wire [31:0] _GEN_23 = _csrData_T_7 ? mideleg_data : _GEN_15; // @[CsrFile.scala 151:31 73:28]
  wire [31:0] _GEN_24 = _csrData_T_7 ? mepc_data : _GEN_16; // @[CsrFile.scala 151:31 74:28]
  wire  _GEN_25 = _csrData_T_7 ? satp_mode : _GEN_17; // @[CsrFile.scala 151:31 75:28]
  wire [21:0] _GEN_26 = _csrData_T_7 ? satp_ppn : _GEN_18; // @[CsrFile.scala 151:31 75:28]
  wire [63:0] _GEN_27 = _csrData_T_7 ? _mcycle_data_T_1 : _GEN_19; // @[CsrFile.scala 148:17 151:31]
  wire [31:0] csrState_mcycle = mcycle_data[31:0]; // @[CsrFile.scala 179:29]
  wire [31:0] csrState_mcycleh = mcycle_data[63:32]; // @[CsrFile.scala 180:30]
  assign io_read_valid = 3'h5 == io_read_op ? _readValid_T : _readValid_T_10; // @[Mux.scala 81:58]
  assign io_read_data = _T_7 ? 32'h0 : _T_97; // @[Lookup.scala 34:39]
  assign io_mepc = mepc_data; // @[CsrFile.scala 173:13]
  assign io_trapVec = {mtvec_base,mtvec_mode}; // @[CsrFile.scala 174:25]
  assign csrState_0_mcycle = csrState_mcycle;
  assign csrState_0_mcycleh = csrState_mcycleh;
  always @(posedge clock) begin
    if (reset) begin // @[CsrFile.scala 69:28]
      mcause_int <= 1'h0; // @[CsrFile.scala 69:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (_csrData_T_3) begin // @[CsrFile.scala 151:31]
        mcause_int <= writeData[31]; // @[CSR.scala 384:11]
      end
    end
    if (reset) begin // @[CsrFile.scala 69:28]
      mcause_code <= 31'h0; // @[CsrFile.scala 69:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (_csrData_T_3) begin // @[CsrFile.scala 151:31]
        mcause_code <= {{27'd0}, writeData[3:0]}; // @[CSR.scala 385:11]
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_sum <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_sum <= writeData[18]; // @[CSR.scala 222:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_mpp <= 2'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_mpp <= writeData[12:11]; // @[CSR.scala 223:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_spp <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_spp <= writeData[8]; // @[CSR.scala 224:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_mpie <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_mpie <= writeData[7]; // @[CSR.scala 225:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_spie <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_spie <= writeData[5]; // @[CSR.scala 226:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_mie <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_mie <= writeData[3]; // @[CSR.scala 227:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_sie <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_sie <= writeData[1]; // @[CSR.scala 228:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 71:28]
      mtvec_base <= 30'h0; // @[CsrFile.scala 71:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          mtvec_base <= _GEN_20;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 71:28]
      mtvec_mode <= 2'h0; // @[CsrFile.scala 71:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          mtvec_mode <= _GEN_21;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 72:28]
      medeleg_data <= 32'h0; // @[CsrFile.scala 72:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          medeleg_data <= _GEN_22;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 73:28]
      mideleg_data <= 32'h0; // @[CsrFile.scala 73:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          mideleg_data <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 74:28]
      mepc_data <= 32'h0; // @[CsrFile.scala 74:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          mepc_data <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 75:28]
      satp_mode <= 1'h0; // @[CsrFile.scala 75:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          satp_mode <= _GEN_25;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 75:28]
      satp_ppn <= 22'h0; // @[CsrFile.scala 75:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          satp_ppn <= _GEN_26;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 77:28]
      mcycle_data <= 64'h0; // @[CsrFile.scala 77:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (_csrData_T_3) begin // @[CsrFile.scala 151:31]
        mcycle_data <= _mcycle_data_T_1; // @[CsrFile.scala 148:17]
      end else if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
        mcycle_data <= _mcycle_data_T_1; // @[CsrFile.scala 148:17]
      end else begin
        mcycle_data <= _GEN_27;
      end
    end else begin
      mcycle_data <= _mcycle_data_T_1; // @[CsrFile.scala 148:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mcause_int = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mcause_code = _RAND_1[30:0];
  _RAND_2 = {1{`RANDOM}};
  mstatus_sum = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  mstatus_mpp = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  mstatus_spp = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  mstatus_mpie = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  mstatus_spie = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  mstatus_mie = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mstatus_sie = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  mtvec_base = _RAND_9[29:0];
  _RAND_10 = {1{`RANDOM}};
  mtvec_mode = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  medeleg_data = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mideleg_data = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mepc_data = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  satp_mode = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  satp_ppn = _RAND_15[21:0];
  _RAND_16 = {2{`RANDOM}};
  mcycle_data = _RAND_16[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSRStage_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [2:0]  io_in_bits_csrOp,
  input  [3:0]  io_in_bits_excpType,
  input  [31:0] io_in_bits_rs1Val,
  input  [31:0] io_in_bits_inst,
  input  [7:0]  io_in_bits_id,
  output        io_out_valid,
  output [4:0]  io_out_bits_rd,
  output [31:0] io_out_bits_data,
  output [31:0] io_out_bits_excpAddr,
  output        io_out_bits_excpValid,
  output [7:0]  io_out_bits_id,
  input         io_flush,
  output [31:0] csrState_mcycle,
  output [31:0] csrState_mcycleh
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  csrFile_clock; // @[CSR.scala 190:25]
  wire  csrFile_reset; // @[CSR.scala 190:25]
  wire [2:0] csrFile_io_read_op; // @[CSR.scala 190:25]
  wire  csrFile_io_read_valid; // @[CSR.scala 190:25]
  wire [11:0] csrFile_io_read_addr; // @[CSR.scala 190:25]
  wire [31:0] csrFile_io_read_data; // @[CSR.scala 190:25]
  wire [2:0] csrFile_io_write_op; // @[CSR.scala 190:25]
  wire [11:0] csrFile_io_write_addr; // @[CSR.scala 190:25]
  wire [31:0] csrFile_io_write_data; // @[CSR.scala 190:25]
  wire [31:0] csrFile_io_mepc; // @[CSR.scala 190:25]
  wire [31:0] csrFile_io_trapVec; // @[CSR.scala 190:25]
  wire [31:0] csrFile_csrState_0_mcycle; // @[CSR.scala 190:25]
  wire [31:0] csrFile_csrState_0_mcycleh; // @[CSR.scala 190:25]
  wire [31:0] immGen_io_inst; // @[CSR.scala 214:24]
  wire [2:0] immGen_io_immSrc; // @[CSR.scala 214:24]
  wire  immGen_io_immSign; // @[CSR.scala 214:24]
  wire [31:0] immGen_io_imm; // @[CSR.scala 214:24]
  reg  s0_full; // @[CSR.scala 206:26]
  reg  s1_full; // @[CSR.scala 240:26]
  wire  s1_ready = ~s1_full | io_out_valid; // @[CSR.scala 250:26]
  wire  s0_fire = s0_full & s1_ready; // @[CSR.scala 207:28]
  wire  s0_ready = ~s0_full | s0_fire; // @[CSR.scala 209:26]
  wire  s0_latch = io_in_valid & s0_ready; // @[CSR.scala 205:32]
  reg [2:0] s0_info_csrOp; // @[Reg.scala 19:16]
  reg [3:0] s0_info_excpType; // @[Reg.scala 19:16]
  reg [31:0] s0_info_rs1Val; // @[Reg.scala 19:16]
  reg [31:0] s0_info_inst; // @[Reg.scala 19:16]
  reg [7:0] s0_info_id; // @[Reg.scala 19:16]
  wire  _GEN_6 = s0_fire & s0_full ? 1'h0 : s0_full; // @[CSR.scala 206:26 212:{35,45}]
  wire  _GEN_7 = s0_latch | _GEN_6; // @[CSR.scala 211:{20,30}]
  wire [11:0] s0_csrAddr = s0_info_inst[31:20]; // @[util.scala 78:36]
  wire  s0_csrWrEn = s0_info_csrOp != 3'h0 & csrFile_io_read_valid; // @[CSR.scala 230:43]
  reg [4:0] s1_rd; // @[Reg.scala 19:16]
  reg [2:0] s1_csrOp; // @[Reg.scala 19:16]
  reg [3:0] s1_excpType; // @[Reg.scala 19:16]
  reg [11:0] s1_csrAddr; // @[Reg.scala 19:16]
  reg  s1_csrWrEn; // @[Reg.scala 19:16]
  reg [31:0] s1_csrWrData; // @[Reg.scala 19:16]
  reg [31:0] s1_csrRdData; // @[Reg.scala 19:16]
  reg [7:0] s1_id; // @[Reg.scala 19:16]
  wire  _GEN_16 = io_out_valid & s1_full ? 1'h0 : s1_full; // @[CSR.scala 240:26 253:{35,45}]
  wire  _GEN_17 = s0_fire | _GEN_16; // @[CSR.scala 252:{20,30}]
  CsrFile csrFile ( // @[CSR.scala 190:25]
    .clock(csrFile_clock),
    .reset(csrFile_reset),
    .io_read_op(csrFile_io_read_op),
    .io_read_valid(csrFile_io_read_valid),
    .io_read_addr(csrFile_io_read_addr),
    .io_read_data(csrFile_io_read_data),
    .io_write_op(csrFile_io_write_op),
    .io_write_addr(csrFile_io_write_addr),
    .io_write_data(csrFile_io_write_data),
    .io_mepc(csrFile_io_mepc),
    .io_trapVec(csrFile_io_trapVec),
    .csrState_0_mcycle(csrFile_csrState_0_mcycle),
    .csrState_0_mcycleh(csrFile_csrState_0_mcycleh)
  );
  ImmGen immGen ( // @[CSR.scala 214:24]
    .io_inst(immGen_io_inst),
    .io_immSrc(immGen_io_immSrc),
    .io_immSign(immGen_io_immSign),
    .io_imm(immGen_io_imm)
  );
  assign io_in_ready = ~s0_full | s0_fire; // @[CSR.scala 209:26]
  assign io_out_valid = s1_full; // @[CSR.scala 266:18]
  assign io_out_bits_rd = s1_rd; // @[CSR.scala 264:20]
  assign io_out_bits_data = s1_csrRdData; // @[CSR.scala 263:22]
  assign io_out_bits_excpAddr = 4'h4 == s1_excpType ? csrFile_io_mepc : csrFile_io_trapVec; // @[Mux.scala 81:58]
  assign io_out_bits_excpValid = s1_excpType != 4'h0; // @[CSR.scala 259:42]
  assign io_out_bits_id = s1_id; // @[CSR.scala 265:20]
  assign csrState_mcycle = csrFile_csrState_0_mcycle;
  assign csrState_mcycleh = csrFile_csrState_0_mcycleh;
  assign csrFile_clock = clock;
  assign csrFile_reset = reset;
  assign csrFile_io_read_op = s0_info_csrOp; // @[CSR.scala 227:24]
  assign csrFile_io_read_addr = s0_info_inst[31:20]; // @[util.scala 78:36]
  assign csrFile_io_write_op = s1_csrWrEn ? s1_csrOp : 3'h1; // @[CSR.scala 257:31]
  assign csrFile_io_write_addr = s1_csrAddr; // @[CSR.scala 255:27]
  assign csrFile_io_write_data = s1_csrWrData; // @[CSR.scala 256:27]
  assign immGen_io_inst = s0_info_inst; // @[CSR.scala 218:20]
  assign immGen_io_immSrc = 3'h5; // @[CSR.scala 216:22]
  assign immGen_io_immSign = 1'h0; // @[CSR.scala 217:23]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 206:26]
      s0_full <= 1'h0; // @[CSR.scala 206:26]
    end else if (io_flush) begin // @[CSR.scala 270:20]
      s0_full <= 1'h0; // @[CSR.scala 271:17]
    end else begin
      s0_full <= _GEN_7;
    end
    if (reset) begin // @[CSR.scala 240:26]
      s1_full <= 1'h0; // @[CSR.scala 240:26]
    end else if (io_flush) begin // @[CSR.scala 270:20]
      s1_full <= 1'h0; // @[CSR.scala 272:17]
    end else begin
      s1_full <= _GEN_17;
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_csrOp <= io_in_bits_csrOp; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_excpType <= io_in_bits_excpType; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_rs1Val <= io_in_bits_rs1Val; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_inst <= io_in_bits_inst; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_info_id <= io_in_bits_id; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rd <= s0_info_inst[11:7]; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_csrOp <= s0_info_csrOp; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_excpType <= s0_info_excpType; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_csrAddr <= s0_csrAddr; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_csrWrEn <= s0_csrWrEn; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_csrWrData <= s0_info_rs1Val; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_csrRdData <= csrFile_io_read_data; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_id <= s0_info_id; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s1_full = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s0_info_csrOp = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  s0_info_excpType = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  s0_info_rs1Val = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  s0_info_inst = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  s0_info_id = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  s1_rd = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  s1_csrOp = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  s1_excpType = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  s1_csrAddr = _RAND_10[11:0];
  _RAND_11 = {1{`RANDOM}};
  s1_csrWrEn = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  s1_csrWrData = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  s1_csrRdData = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  s1_id = _RAND_14[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EdgeDetect(
  input   clock,
  input   io_in,
  output  io_change
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  prev; // @[Core_1.scala 27:23]
  assign io_change = prev & ~io_in; // @[Core_1.scala 31:27]
  always @(posedge clock) begin
    prev <= io_in; // @[Core_1.scala 27:23]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prev = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_5(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits = empty ? io_enq_bits : ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decoder_1(
  input  [31:0] io_inst,
  output [3:0]  io_out_brType,
  output [2:0]  io_out_wbType,
  output [4:0]  io_out_lsuOp,
  output [4:0]  io_out_aluOp,
  output [3:0]  io_out_opr1,
  output [3:0]  io_out_opr2,
  output [2:0]  io_out_immSrc,
  output        io_out_immSign,
  output [2:0]  io_out_csrOp,
  output [3:0]  io_out_excpType
);
  wire [31:0] _decodeSigs_T = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_1 = 32'h3 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_3 = 32'h1003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_5 = 32'h2003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_7 = 32'h4003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_9 = 32'h5003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_11 = 32'h13 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [31:0] _decodeSigs_T_12 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_13 = 32'h1013 == _decodeSigs_T_12; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_15 = 32'h2013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_17 = 32'h3013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_19 = 32'h4013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_21 = 32'h5013 == _decodeSigs_T_12; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_23 = 32'h40005013 == _decodeSigs_T_12; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_25 = 32'h6013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_27 = 32'h7013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [31:0] _decodeSigs_T_28 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_29 = 32'h17 == _decodeSigs_T_28; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_31 = 32'h23 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_33 = 32'h1023 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_35 = 32'h2023 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [31:0] _decodeSigs_T_36 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_37 = 32'h33 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_39 = 32'h40000033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_41 = 32'h1033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_43 = 32'h2033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_45 = 32'h3033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_47 = 32'h4033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_49 = 32'h5033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_51 = 32'h40005033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_53 = 32'h6033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_55 = 32'h7033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_57 = 32'h37 == _decodeSigs_T_28; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_59 = 32'h63 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_61 = 32'h1063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_63 = 32'h4063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_65 = 32'h5063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_67 = 32'h6063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_69 = 32'h7063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_71 = 32'h67 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_73 = 32'h6f == _decodeSigs_T_28; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_75 = 32'hf == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_77 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_79 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_81 = 32'h30200073 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_83 = 32'h10200073 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_85 = 32'h1073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_87 = 32'h2073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_89 = 32'h3073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_91 = 32'h5073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_93 = 32'h6073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_95 = 32'h7073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [3:0] _decodeSigs_T_107 = _decodeSigs_T_73 ? 4'h1 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_108 = _decodeSigs_T_71 ? 4'h2 : _decodeSigs_T_107; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_109 = _decodeSigs_T_69 ? 4'h8 : _decodeSigs_T_108; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_110 = _decodeSigs_T_67 ? 4'h7 : _decodeSigs_T_109; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_111 = _decodeSigs_T_65 ? 4'h5 : _decodeSigs_T_110; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_112 = _decodeSigs_T_63 ? 4'h6 : _decodeSigs_T_111; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_113 = _decodeSigs_T_61 ? 4'h4 : _decodeSigs_T_112; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_114 = _decodeSigs_T_59 ? 4'h3 : _decodeSigs_T_113; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_115 = _decodeSigs_T_57 ? 4'h0 : _decodeSigs_T_114; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_116 = _decodeSigs_T_55 ? 4'h0 : _decodeSigs_T_115; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_117 = _decodeSigs_T_53 ? 4'h0 : _decodeSigs_T_116; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_118 = _decodeSigs_T_51 ? 4'h0 : _decodeSigs_T_117; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_119 = _decodeSigs_T_49 ? 4'h0 : _decodeSigs_T_118; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_120 = _decodeSigs_T_47 ? 4'h0 : _decodeSigs_T_119; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_121 = _decodeSigs_T_45 ? 4'h0 : _decodeSigs_T_120; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_122 = _decodeSigs_T_43 ? 4'h0 : _decodeSigs_T_121; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_123 = _decodeSigs_T_41 ? 4'h0 : _decodeSigs_T_122; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_124 = _decodeSigs_T_39 ? 4'h0 : _decodeSigs_T_123; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_125 = _decodeSigs_T_37 ? 4'h0 : _decodeSigs_T_124; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_126 = _decodeSigs_T_35 ? 4'h0 : _decodeSigs_T_125; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_127 = _decodeSigs_T_33 ? 4'h0 : _decodeSigs_T_126; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_128 = _decodeSigs_T_31 ? 4'h0 : _decodeSigs_T_127; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_129 = _decodeSigs_T_29 ? 4'h0 : _decodeSigs_T_128; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_130 = _decodeSigs_T_27 ? 4'h0 : _decodeSigs_T_129; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_131 = _decodeSigs_T_25 ? 4'h0 : _decodeSigs_T_130; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_132 = _decodeSigs_T_23 ? 4'h0 : _decodeSigs_T_131; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_133 = _decodeSigs_T_21 ? 4'h0 : _decodeSigs_T_132; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_134 = _decodeSigs_T_19 ? 4'h0 : _decodeSigs_T_133; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_135 = _decodeSigs_T_17 ? 4'h0 : _decodeSigs_T_134; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_136 = _decodeSigs_T_15 ? 4'h0 : _decodeSigs_T_135; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_137 = _decodeSigs_T_13 ? 4'h0 : _decodeSigs_T_136; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_138 = _decodeSigs_T_11 ? 4'h0 : _decodeSigs_T_137; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_139 = _decodeSigs_T_9 ? 4'h0 : _decodeSigs_T_138; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_140 = _decodeSigs_T_7 ? 4'h0 : _decodeSigs_T_139; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_141 = _decodeSigs_T_5 ? 4'h0 : _decodeSigs_T_140; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_142 = _decodeSigs_T_3 ? 4'h0 : _decodeSigs_T_141; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_143 = _decodeSigs_T_95 ? 3'h4 : 3'h1; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_144 = _decodeSigs_T_93 ? 3'h4 : _decodeSigs_T_143; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_145 = _decodeSigs_T_91 ? 3'h4 : _decodeSigs_T_144; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_146 = _decodeSigs_T_89 ? 3'h4 : _decodeSigs_T_145; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_147 = _decodeSigs_T_87 ? 3'h4 : _decodeSigs_T_146; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_148 = _decodeSigs_T_85 ? 3'h4 : _decodeSigs_T_147; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_149 = _decodeSigs_T_83 ? 3'h1 : _decodeSigs_T_148; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_150 = _decodeSigs_T_81 ? 3'h1 : _decodeSigs_T_149; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_151 = _decodeSigs_T_79 ? 3'h1 : _decodeSigs_T_150; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_152 = _decodeSigs_T_77 ? 3'h1 : _decodeSigs_T_151; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_153 = _decodeSigs_T_75 ? 3'h1 : _decodeSigs_T_152; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_154 = _decodeSigs_T_73 ? 3'h3 : _decodeSigs_T_153; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_155 = _decodeSigs_T_71 ? 3'h3 : _decodeSigs_T_154; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_156 = _decodeSigs_T_69 ? 3'h1 : _decodeSigs_T_155; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_157 = _decodeSigs_T_67 ? 3'h1 : _decodeSigs_T_156; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_158 = _decodeSigs_T_65 ? 3'h1 : _decodeSigs_T_157; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_159 = _decodeSigs_T_63 ? 3'h1 : _decodeSigs_T_158; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_160 = _decodeSigs_T_61 ? 3'h1 : _decodeSigs_T_159; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_161 = _decodeSigs_T_59 ? 3'h1 : _decodeSigs_T_160; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_162 = _decodeSigs_T_57 ? 3'h1 : _decodeSigs_T_161; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_163 = _decodeSigs_T_55 ? 3'h1 : _decodeSigs_T_162; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_164 = _decodeSigs_T_53 ? 3'h1 : _decodeSigs_T_163; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_165 = _decodeSigs_T_51 ? 3'h1 : _decodeSigs_T_164; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_166 = _decodeSigs_T_49 ? 3'h1 : _decodeSigs_T_165; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_167 = _decodeSigs_T_47 ? 3'h1 : _decodeSigs_T_166; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_168 = _decodeSigs_T_45 ? 3'h1 : _decodeSigs_T_167; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_169 = _decodeSigs_T_43 ? 3'h1 : _decodeSigs_T_168; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_170 = _decodeSigs_T_41 ? 3'h1 : _decodeSigs_T_169; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_171 = _decodeSigs_T_39 ? 3'h1 : _decodeSigs_T_170; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_172 = _decodeSigs_T_37 ? 3'h1 : _decodeSigs_T_171; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_173 = _decodeSigs_T_35 ? 3'h0 : _decodeSigs_T_172; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_174 = _decodeSigs_T_33 ? 3'h0 : _decodeSigs_T_173; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_175 = _decodeSigs_T_31 ? 3'h0 : _decodeSigs_T_174; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_176 = _decodeSigs_T_29 ? 3'h1 : _decodeSigs_T_175; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_177 = _decodeSigs_T_27 ? 3'h1 : _decodeSigs_T_176; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_178 = _decodeSigs_T_25 ? 3'h1 : _decodeSigs_T_177; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_179 = _decodeSigs_T_23 ? 3'h1 : _decodeSigs_T_178; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_180 = _decodeSigs_T_21 ? 3'h1 : _decodeSigs_T_179; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_181 = _decodeSigs_T_19 ? 3'h1 : _decodeSigs_T_180; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_182 = _decodeSigs_T_17 ? 3'h1 : _decodeSigs_T_181; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_183 = _decodeSigs_T_15 ? 3'h1 : _decodeSigs_T_182; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_184 = _decodeSigs_T_13 ? 3'h1 : _decodeSigs_T_183; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_185 = _decodeSigs_T_11 ? 3'h1 : _decodeSigs_T_184; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_186 = _decodeSigs_T_9 ? 3'h2 : _decodeSigs_T_185; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_187 = _decodeSigs_T_7 ? 3'h2 : _decodeSigs_T_186; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_188 = _decodeSigs_T_5 ? 3'h2 : _decodeSigs_T_187; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_189 = _decodeSigs_T_3 ? 3'h2 : _decodeSigs_T_188; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_200 = _decodeSigs_T_75 ? 5'h14 : 5'h0; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_201 = _decodeSigs_T_73 ? 5'h0 : _decodeSigs_T_200; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_202 = _decodeSigs_T_71 ? 5'h0 : _decodeSigs_T_201; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_203 = _decodeSigs_T_69 ? 5'h0 : _decodeSigs_T_202; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_204 = _decodeSigs_T_67 ? 5'h0 : _decodeSigs_T_203; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_205 = _decodeSigs_T_65 ? 5'h0 : _decodeSigs_T_204; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_206 = _decodeSigs_T_63 ? 5'h0 : _decodeSigs_T_205; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_207 = _decodeSigs_T_61 ? 5'h0 : _decodeSigs_T_206; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_208 = _decodeSigs_T_59 ? 5'h0 : _decodeSigs_T_207; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_209 = _decodeSigs_T_57 ? 5'h0 : _decodeSigs_T_208; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_210 = _decodeSigs_T_55 ? 5'h0 : _decodeSigs_T_209; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_211 = _decodeSigs_T_53 ? 5'h0 : _decodeSigs_T_210; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_212 = _decodeSigs_T_51 ? 5'h0 : _decodeSigs_T_211; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_213 = _decodeSigs_T_49 ? 5'h0 : _decodeSigs_T_212; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_214 = _decodeSigs_T_47 ? 5'h0 : _decodeSigs_T_213; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_215 = _decodeSigs_T_45 ? 5'h0 : _decodeSigs_T_214; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_216 = _decodeSigs_T_43 ? 5'h0 : _decodeSigs_T_215; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_217 = _decodeSigs_T_41 ? 5'h0 : _decodeSigs_T_216; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_218 = _decodeSigs_T_39 ? 5'h0 : _decodeSigs_T_217; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_219 = _decodeSigs_T_37 ? 5'h0 : _decodeSigs_T_218; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_220 = _decodeSigs_T_35 ? 5'h8 : _decodeSigs_T_219; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_221 = _decodeSigs_T_33 ? 5'h7 : _decodeSigs_T_220; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_222 = _decodeSigs_T_31 ? 5'h6 : _decodeSigs_T_221; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_223 = _decodeSigs_T_29 ? 5'h0 : _decodeSigs_T_222; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_224 = _decodeSigs_T_27 ? 5'h0 : _decodeSigs_T_223; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_225 = _decodeSigs_T_25 ? 5'h0 : _decodeSigs_T_224; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_226 = _decodeSigs_T_23 ? 5'h0 : _decodeSigs_T_225; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_227 = _decodeSigs_T_21 ? 5'h0 : _decodeSigs_T_226; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_228 = _decodeSigs_T_19 ? 5'h0 : _decodeSigs_T_227; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_229 = _decodeSigs_T_17 ? 5'h0 : _decodeSigs_T_228; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_230 = _decodeSigs_T_15 ? 5'h0 : _decodeSigs_T_229; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_231 = _decodeSigs_T_13 ? 5'h0 : _decodeSigs_T_230; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_232 = _decodeSigs_T_11 ? 5'h0 : _decodeSigs_T_231; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_233 = _decodeSigs_T_9 ? 5'h5 : _decodeSigs_T_232; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_234 = _decodeSigs_T_7 ? 5'h4 : _decodeSigs_T_233; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_235 = _decodeSigs_T_5 ? 5'h3 : _decodeSigs_T_234; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_236 = _decodeSigs_T_3 ? 5'h2 : _decodeSigs_T_235; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_256 = _decodeSigs_T_57 ? 5'h0 : 5'h11; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_257 = _decodeSigs_T_55 ? 5'h2 : _decodeSigs_T_256; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_258 = _decodeSigs_T_53 ? 5'h3 : _decodeSigs_T_257; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_259 = _decodeSigs_T_51 ? 5'hc : _decodeSigs_T_258; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_260 = _decodeSigs_T_49 ? 5'hb : _decodeSigs_T_259; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_261 = _decodeSigs_T_47 ? 5'h4 : _decodeSigs_T_260; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_262 = _decodeSigs_T_45 ? 5'h9 : _decodeSigs_T_261; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_263 = _decodeSigs_T_43 ? 5'h8 : _decodeSigs_T_262; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_264 = _decodeSigs_T_41 ? 5'ha : _decodeSigs_T_263; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_265 = _decodeSigs_T_39 ? 5'h1 : _decodeSigs_T_264; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_266 = _decodeSigs_T_37 ? 5'h0 : _decodeSigs_T_265; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_267 = _decodeSigs_T_35 ? 5'h11 : _decodeSigs_T_266; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_268 = _decodeSigs_T_33 ? 5'h11 : _decodeSigs_T_267; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_269 = _decodeSigs_T_31 ? 5'h11 : _decodeSigs_T_268; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_270 = _decodeSigs_T_29 ? 5'h0 : _decodeSigs_T_269; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_271 = _decodeSigs_T_27 ? 5'h2 : _decodeSigs_T_270; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_272 = _decodeSigs_T_25 ? 5'h3 : _decodeSigs_T_271; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_273 = _decodeSigs_T_23 ? 5'hc : _decodeSigs_T_272; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_274 = _decodeSigs_T_21 ? 5'hb : _decodeSigs_T_273; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_275 = _decodeSigs_T_19 ? 5'h4 : _decodeSigs_T_274; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_276 = _decodeSigs_T_17 ? 5'h9 : _decodeSigs_T_275; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_277 = _decodeSigs_T_15 ? 5'h8 : _decodeSigs_T_276; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_278 = _decodeSigs_T_13 ? 5'ha : _decodeSigs_T_277; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_279 = _decodeSigs_T_11 ? 5'h0 : _decodeSigs_T_278; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_280 = _decodeSigs_T_9 ? 5'h11 : _decodeSigs_T_279; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_281 = _decodeSigs_T_7 ? 5'h11 : _decodeSigs_T_280; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_282 = _decodeSigs_T_5 ? 5'h11 : _decodeSigs_T_281; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_283 = _decodeSigs_T_3 ? 5'h11 : _decodeSigs_T_282; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_284 = _decodeSigs_T_95 ? 4'h6 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_285 = _decodeSigs_T_93 ? 4'h6 : _decodeSigs_T_284; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_286 = _decodeSigs_T_91 ? 4'h6 : _decodeSigs_T_285; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_287 = _decodeSigs_T_89 ? 4'h1 : _decodeSigs_T_286; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_288 = _decodeSigs_T_87 ? 4'h1 : _decodeSigs_T_287; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_289 = _decodeSigs_T_85 ? 4'h1 : _decodeSigs_T_288; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_290 = _decodeSigs_T_83 ? 4'h0 : _decodeSigs_T_289; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_291 = _decodeSigs_T_81 ? 4'h0 : _decodeSigs_T_290; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_292 = _decodeSigs_T_79 ? 4'h0 : _decodeSigs_T_291; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_293 = _decodeSigs_T_77 ? 4'h0 : _decodeSigs_T_292; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_294 = _decodeSigs_T_75 ? 4'h0 : _decodeSigs_T_293; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_295 = _decodeSigs_T_73 ? 4'h7 : _decodeSigs_T_294; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_296 = _decodeSigs_T_71 ? 4'h1 : _decodeSigs_T_295; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_297 = _decodeSigs_T_69 ? 4'h1 : _decodeSigs_T_296; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_298 = _decodeSigs_T_67 ? 4'h1 : _decodeSigs_T_297; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_299 = _decodeSigs_T_65 ? 4'h1 : _decodeSigs_T_298; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_300 = _decodeSigs_T_63 ? 4'h1 : _decodeSigs_T_299; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_301 = _decodeSigs_T_61 ? 4'h1 : _decodeSigs_T_300; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_302 = _decodeSigs_T_59 ? 4'h1 : _decodeSigs_T_301; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_303 = _decodeSigs_T_57 ? 4'h0 : _decodeSigs_T_302; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_304 = _decodeSigs_T_55 ? 4'h1 : _decodeSigs_T_303; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_305 = _decodeSigs_T_53 ? 4'h1 : _decodeSigs_T_304; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_306 = _decodeSigs_T_51 ? 4'h1 : _decodeSigs_T_305; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_307 = _decodeSigs_T_49 ? 4'h1 : _decodeSigs_T_306; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_308 = _decodeSigs_T_47 ? 4'h1 : _decodeSigs_T_307; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_309 = _decodeSigs_T_45 ? 4'h1 : _decodeSigs_T_308; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_310 = _decodeSigs_T_43 ? 4'h1 : _decodeSigs_T_309; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_311 = _decodeSigs_T_41 ? 4'h1 : _decodeSigs_T_310; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_312 = _decodeSigs_T_39 ? 4'h1 : _decodeSigs_T_311; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_313 = _decodeSigs_T_37 ? 4'h1 : _decodeSigs_T_312; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_314 = _decodeSigs_T_35 ? 4'h1 : _decodeSigs_T_313; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_315 = _decodeSigs_T_33 ? 4'h1 : _decodeSigs_T_314; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_316 = _decodeSigs_T_31 ? 4'h1 : _decodeSigs_T_315; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_317 = _decodeSigs_T_29 ? 4'h7 : _decodeSigs_T_316; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_318 = _decodeSigs_T_27 ? 4'h1 : _decodeSigs_T_317; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_319 = _decodeSigs_T_25 ? 4'h1 : _decodeSigs_T_318; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_320 = _decodeSigs_T_23 ? 4'h1 : _decodeSigs_T_319; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_321 = _decodeSigs_T_21 ? 4'h1 : _decodeSigs_T_320; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_322 = _decodeSigs_T_19 ? 4'h1 : _decodeSigs_T_321; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_323 = _decodeSigs_T_17 ? 4'h1 : _decodeSigs_T_322; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_324 = _decodeSigs_T_15 ? 4'h1 : _decodeSigs_T_323; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_325 = _decodeSigs_T_13 ? 4'h1 : _decodeSigs_T_324; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_326 = _decodeSigs_T_11 ? 4'h1 : _decodeSigs_T_325; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_327 = _decodeSigs_T_9 ? 4'h1 : _decodeSigs_T_326; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_328 = _decodeSigs_T_7 ? 4'h1 : _decodeSigs_T_327; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_329 = _decodeSigs_T_5 ? 4'h1 : _decodeSigs_T_328; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_330 = _decodeSigs_T_3 ? 4'h1 : _decodeSigs_T_329; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_342 = _decodeSigs_T_73 ? 4'h3 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_343 = _decodeSigs_T_71 ? 4'h3 : _decodeSigs_T_342; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_344 = _decodeSigs_T_69 ? 4'h2 : _decodeSigs_T_343; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_345 = _decodeSigs_T_67 ? 4'h2 : _decodeSigs_T_344; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_346 = _decodeSigs_T_65 ? 4'h2 : _decodeSigs_T_345; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_347 = _decodeSigs_T_63 ? 4'h2 : _decodeSigs_T_346; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_348 = _decodeSigs_T_61 ? 4'h2 : _decodeSigs_T_347; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_349 = _decodeSigs_T_59 ? 4'h2 : _decodeSigs_T_348; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_350 = _decodeSigs_T_57 ? 4'h3 : _decodeSigs_T_349; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_351 = _decodeSigs_T_55 ? 4'h2 : _decodeSigs_T_350; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_352 = _decodeSigs_T_53 ? 4'h2 : _decodeSigs_T_351; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_353 = _decodeSigs_T_51 ? 4'h2 : _decodeSigs_T_352; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_354 = _decodeSigs_T_49 ? 4'h2 : _decodeSigs_T_353; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_355 = _decodeSigs_T_47 ? 4'h2 : _decodeSigs_T_354; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_356 = _decodeSigs_T_45 ? 4'h2 : _decodeSigs_T_355; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_357 = _decodeSigs_T_43 ? 4'h2 : _decodeSigs_T_356; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_358 = _decodeSigs_T_41 ? 4'h2 : _decodeSigs_T_357; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_359 = _decodeSigs_T_39 ? 4'h2 : _decodeSigs_T_358; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_360 = _decodeSigs_T_37 ? 4'h2 : _decodeSigs_T_359; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_361 = _decodeSigs_T_35 ? 4'h2 : _decodeSigs_T_360; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_362 = _decodeSigs_T_33 ? 4'h2 : _decodeSigs_T_361; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_363 = _decodeSigs_T_31 ? 4'h2 : _decodeSigs_T_362; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_364 = _decodeSigs_T_29 ? 4'h3 : _decodeSigs_T_363; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_365 = _decodeSigs_T_27 ? 4'h3 : _decodeSigs_T_364; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_366 = _decodeSigs_T_25 ? 4'h3 : _decodeSigs_T_365; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_367 = _decodeSigs_T_23 ? 4'h3 : _decodeSigs_T_366; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_368 = _decodeSigs_T_21 ? 4'h3 : _decodeSigs_T_367; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_369 = _decodeSigs_T_19 ? 4'h3 : _decodeSigs_T_368; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_370 = _decodeSigs_T_17 ? 4'h3 : _decodeSigs_T_369; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_371 = _decodeSigs_T_15 ? 4'h3 : _decodeSigs_T_370; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_372 = _decodeSigs_T_13 ? 4'h3 : _decodeSigs_T_371; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_373 = _decodeSigs_T_11 ? 4'h3 : _decodeSigs_T_372; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_374 = _decodeSigs_T_9 ? 4'h0 : _decodeSigs_T_373; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_375 = _decodeSigs_T_7 ? 4'h0 : _decodeSigs_T_374; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_376 = _decodeSigs_T_5 ? 4'h0 : _decodeSigs_T_375; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_377 = _decodeSigs_T_3 ? 4'h0 : _decodeSigs_T_376; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_378 = _decodeSigs_T_95 ? 3'h5 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_379 = _decodeSigs_T_93 ? 3'h5 : _decodeSigs_T_378; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_380 = _decodeSigs_T_91 ? 3'h5 : _decodeSigs_T_379; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_381 = _decodeSigs_T_89 ? 3'h0 : _decodeSigs_T_380; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_382 = _decodeSigs_T_87 ? 3'h0 : _decodeSigs_T_381; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_383 = _decodeSigs_T_85 ? 3'h0 : _decodeSigs_T_382; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_384 = _decodeSigs_T_83 ? 3'h0 : _decodeSigs_T_383; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_385 = _decodeSigs_T_81 ? 3'h0 : _decodeSigs_T_384; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_386 = _decodeSigs_T_79 ? 3'h0 : _decodeSigs_T_385; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_387 = _decodeSigs_T_77 ? 3'h0 : _decodeSigs_T_386; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_388 = _decodeSigs_T_75 ? 3'h0 : _decodeSigs_T_387; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_389 = _decodeSigs_T_73 ? 3'h4 : _decodeSigs_T_388; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_390 = _decodeSigs_T_71 ? 3'h0 : _decodeSigs_T_389; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_391 = _decodeSigs_T_69 ? 3'h2 : _decodeSigs_T_390; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_392 = _decodeSigs_T_67 ? 3'h2 : _decodeSigs_T_391; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_393 = _decodeSigs_T_65 ? 3'h2 : _decodeSigs_T_392; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_394 = _decodeSigs_T_63 ? 3'h2 : _decodeSigs_T_393; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_395 = _decodeSigs_T_61 ? 3'h2 : _decodeSigs_T_394; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_396 = _decodeSigs_T_59 ? 3'h2 : _decodeSigs_T_395; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_397 = _decodeSigs_T_57 ? 3'h3 : _decodeSigs_T_396; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_398 = _decodeSigs_T_55 ? 3'h0 : _decodeSigs_T_397; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_399 = _decodeSigs_T_53 ? 3'h0 : _decodeSigs_T_398; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_400 = _decodeSigs_T_51 ? 3'h0 : _decodeSigs_T_399; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_401 = _decodeSigs_T_49 ? 3'h0 : _decodeSigs_T_400; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_402 = _decodeSigs_T_47 ? 3'h0 : _decodeSigs_T_401; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_403 = _decodeSigs_T_45 ? 3'h0 : _decodeSigs_T_402; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_404 = _decodeSigs_T_43 ? 3'h0 : _decodeSigs_T_403; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_405 = _decodeSigs_T_41 ? 3'h0 : _decodeSigs_T_404; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_406 = _decodeSigs_T_39 ? 3'h0 : _decodeSigs_T_405; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_407 = _decodeSigs_T_37 ? 3'h0 : _decodeSigs_T_406; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_408 = _decodeSigs_T_35 ? 3'h1 : _decodeSigs_T_407; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_409 = _decodeSigs_T_33 ? 3'h1 : _decodeSigs_T_408; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_410 = _decodeSigs_T_31 ? 3'h1 : _decodeSigs_T_409; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_411 = _decodeSigs_T_29 ? 3'h3 : _decodeSigs_T_410; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_412 = _decodeSigs_T_27 ? 3'h0 : _decodeSigs_T_411; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_413 = _decodeSigs_T_25 ? 3'h0 : _decodeSigs_T_412; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_414 = _decodeSigs_T_23 ? 3'h0 : _decodeSigs_T_413; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_415 = _decodeSigs_T_21 ? 3'h0 : _decodeSigs_T_414; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_416 = _decodeSigs_T_19 ? 3'h0 : _decodeSigs_T_415; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_417 = _decodeSigs_T_17 ? 3'h0 : _decodeSigs_T_416; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_418 = _decodeSigs_T_15 ? 3'h0 : _decodeSigs_T_417; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_419 = _decodeSigs_T_13 ? 3'h0 : _decodeSigs_T_418; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_420 = _decodeSigs_T_11 ? 3'h0 : _decodeSigs_T_419; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_421 = _decodeSigs_T_9 ? 3'h0 : _decodeSigs_T_420; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_422 = _decodeSigs_T_7 ? 3'h0 : _decodeSigs_T_421; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_423 = _decodeSigs_T_5 ? 3'h0 : _decodeSigs_T_422; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_424 = _decodeSigs_T_3 ? 3'h0 : _decodeSigs_T_423; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_425 = _decodeSigs_T_95 ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_426 = _decodeSigs_T_93 ? 1'h0 : _decodeSigs_T_425; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_427 = _decodeSigs_T_91 ? 1'h0 : _decodeSigs_T_426; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_428 = _decodeSigs_T_89 ? 1'h0 : _decodeSigs_T_427; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_429 = _decodeSigs_T_87 ? 1'h0 : _decodeSigs_T_428; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_430 = _decodeSigs_T_85 ? 1'h0 : _decodeSigs_T_429; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_431 = _decodeSigs_T_83 ? 1'h0 : _decodeSigs_T_430; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_432 = _decodeSigs_T_81 ? 1'h0 : _decodeSigs_T_431; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_433 = _decodeSigs_T_79 ? 1'h0 : _decodeSigs_T_432; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_434 = _decodeSigs_T_77 ? 1'h0 : _decodeSigs_T_433; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_444 = _decodeSigs_T_57 ? 1'h0 : _decodeSigs_T_59 | (_decodeSigs_T_61 | (_decodeSigs_T_63 | (
    _decodeSigs_T_65 | (_decodeSigs_T_67 | (_decodeSigs_T_69 | (_decodeSigs_T_71 | (_decodeSigs_T_73 | (_decodeSigs_T_75
     | _decodeSigs_T_434)))))))); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_445 = _decodeSigs_T_55 ? 1'h0 : _decodeSigs_T_444; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_446 = _decodeSigs_T_53 ? 1'h0 : _decodeSigs_T_445; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_447 = _decodeSigs_T_51 ? 1'h0 : _decodeSigs_T_446; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_448 = _decodeSigs_T_49 ? 1'h0 : _decodeSigs_T_447; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_449 = _decodeSigs_T_47 ? 1'h0 : _decodeSigs_T_448; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_450 = _decodeSigs_T_45 ? 1'h0 : _decodeSigs_T_449; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_451 = _decodeSigs_T_43 ? 1'h0 : _decodeSigs_T_450; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_452 = _decodeSigs_T_41 ? 1'h0 : _decodeSigs_T_451; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_453 = _decodeSigs_T_39 ? 1'h0 : _decodeSigs_T_452; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_454 = _decodeSigs_T_37 ? 1'h0 : _decodeSigs_T_453; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_458 = _decodeSigs_T_29 ? 1'h0 : _decodeSigs_T_31 | (_decodeSigs_T_33 | (_decodeSigs_T_35 |
    _decodeSigs_T_454)); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_462 = _decodeSigs_T_21 ? 1'h0 : _decodeSigs_T_23 | (_decodeSigs_T_25 | (_decodeSigs_T_27 |
    _decodeSigs_T_458)); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_466 = _decodeSigs_T_13 ? 1'h0 : _decodeSigs_T_15 | (_decodeSigs_T_17 | (_decodeSigs_T_19 |
    _decodeSigs_T_462)); // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_473 = _decodeSigs_T_93 ? 3'h4 : _decodeSigs_T_378; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_474 = _decodeSigs_T_91 ? 3'h3 : _decodeSigs_T_473; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_475 = _decodeSigs_T_89 ? 3'h5 : _decodeSigs_T_474; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_476 = _decodeSigs_T_87 ? 3'h4 : _decodeSigs_T_475; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_477 = _decodeSigs_T_85 ? 3'h3 : _decodeSigs_T_476; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_478 = _decodeSigs_T_83 ? 3'h0 : _decodeSigs_T_477; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_479 = _decodeSigs_T_81 ? 3'h0 : _decodeSigs_T_478; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_480 = _decodeSigs_T_79 ? 3'h0 : _decodeSigs_T_479; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_481 = _decodeSigs_T_77 ? 3'h0 : _decodeSigs_T_480; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_482 = _decodeSigs_T_75 ? 3'h0 : _decodeSigs_T_481; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_483 = _decodeSigs_T_73 ? 3'h0 : _decodeSigs_T_482; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_484 = _decodeSigs_T_71 ? 3'h0 : _decodeSigs_T_483; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_485 = _decodeSigs_T_69 ? 3'h0 : _decodeSigs_T_484; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_486 = _decodeSigs_T_67 ? 3'h0 : _decodeSigs_T_485; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_487 = _decodeSigs_T_65 ? 3'h0 : _decodeSigs_T_486; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_488 = _decodeSigs_T_63 ? 3'h0 : _decodeSigs_T_487; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_489 = _decodeSigs_T_61 ? 3'h0 : _decodeSigs_T_488; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_490 = _decodeSigs_T_59 ? 3'h0 : _decodeSigs_T_489; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_491 = _decodeSigs_T_57 ? 3'h0 : _decodeSigs_T_490; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_492 = _decodeSigs_T_55 ? 3'h0 : _decodeSigs_T_491; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_493 = _decodeSigs_T_53 ? 3'h0 : _decodeSigs_T_492; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_494 = _decodeSigs_T_51 ? 3'h0 : _decodeSigs_T_493; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_495 = _decodeSigs_T_49 ? 3'h0 : _decodeSigs_T_494; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_496 = _decodeSigs_T_47 ? 3'h0 : _decodeSigs_T_495; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_497 = _decodeSigs_T_45 ? 3'h0 : _decodeSigs_T_496; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_498 = _decodeSigs_T_43 ? 3'h0 : _decodeSigs_T_497; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_499 = _decodeSigs_T_41 ? 3'h0 : _decodeSigs_T_498; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_500 = _decodeSigs_T_39 ? 3'h0 : _decodeSigs_T_499; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_501 = _decodeSigs_T_37 ? 3'h0 : _decodeSigs_T_500; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_502 = _decodeSigs_T_35 ? 3'h0 : _decodeSigs_T_501; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_503 = _decodeSigs_T_33 ? 3'h0 : _decodeSigs_T_502; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_504 = _decodeSigs_T_31 ? 3'h0 : _decodeSigs_T_503; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_505 = _decodeSigs_T_29 ? 3'h0 : _decodeSigs_T_504; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_506 = _decodeSigs_T_27 ? 3'h0 : _decodeSigs_T_505; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_507 = _decodeSigs_T_25 ? 3'h0 : _decodeSigs_T_506; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_508 = _decodeSigs_T_23 ? 3'h0 : _decodeSigs_T_507; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_509 = _decodeSigs_T_21 ? 3'h0 : _decodeSigs_T_508; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_510 = _decodeSigs_T_19 ? 3'h0 : _decodeSigs_T_509; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_511 = _decodeSigs_T_17 ? 3'h0 : _decodeSigs_T_510; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_512 = _decodeSigs_T_15 ? 3'h0 : _decodeSigs_T_511; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_513 = _decodeSigs_T_13 ? 3'h0 : _decodeSigs_T_512; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_514 = _decodeSigs_T_11 ? 3'h0 : _decodeSigs_T_513; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_515 = _decodeSigs_T_9 ? 3'h0 : _decodeSigs_T_514; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_516 = _decodeSigs_T_7 ? 3'h0 : _decodeSigs_T_515; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_517 = _decodeSigs_T_5 ? 3'h0 : _decodeSigs_T_516; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_518 = _decodeSigs_T_3 ? 3'h0 : _decodeSigs_T_517; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_519 = _decodeSigs_T_95 ? 4'h0 : 4'h5; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_520 = _decodeSigs_T_93 ? 4'h0 : _decodeSigs_T_519; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_521 = _decodeSigs_T_91 ? 4'h0 : _decodeSigs_T_520; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_522 = _decodeSigs_T_89 ? 4'h0 : _decodeSigs_T_521; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_523 = _decodeSigs_T_87 ? 4'h0 : _decodeSigs_T_522; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_524 = _decodeSigs_T_85 ? 4'h0 : _decodeSigs_T_523; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_525 = _decodeSigs_T_83 ? 4'h3 : _decodeSigs_T_524; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_526 = _decodeSigs_T_81 ? 4'h4 : _decodeSigs_T_525; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_527 = _decodeSigs_T_79 ? 4'h2 : _decodeSigs_T_526; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_528 = _decodeSigs_T_77 ? 4'h1 : _decodeSigs_T_527; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_529 = _decodeSigs_T_75 ? 4'h0 : _decodeSigs_T_528; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_530 = _decodeSigs_T_73 ? 4'h0 : _decodeSigs_T_529; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_531 = _decodeSigs_T_71 ? 4'h0 : _decodeSigs_T_530; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_532 = _decodeSigs_T_69 ? 4'h0 : _decodeSigs_T_531; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_533 = _decodeSigs_T_67 ? 4'h0 : _decodeSigs_T_532; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_534 = _decodeSigs_T_65 ? 4'h0 : _decodeSigs_T_533; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_535 = _decodeSigs_T_63 ? 4'h0 : _decodeSigs_T_534; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_536 = _decodeSigs_T_61 ? 4'h0 : _decodeSigs_T_535; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_537 = _decodeSigs_T_59 ? 4'h0 : _decodeSigs_T_536; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_538 = _decodeSigs_T_57 ? 4'h0 : _decodeSigs_T_537; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_539 = _decodeSigs_T_55 ? 4'h0 : _decodeSigs_T_538; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_540 = _decodeSigs_T_53 ? 4'h0 : _decodeSigs_T_539; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_541 = _decodeSigs_T_51 ? 4'h0 : _decodeSigs_T_540; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_542 = _decodeSigs_T_49 ? 4'h0 : _decodeSigs_T_541; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_543 = _decodeSigs_T_47 ? 4'h0 : _decodeSigs_T_542; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_544 = _decodeSigs_T_45 ? 4'h0 : _decodeSigs_T_543; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_545 = _decodeSigs_T_43 ? 4'h0 : _decodeSigs_T_544; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_546 = _decodeSigs_T_41 ? 4'h0 : _decodeSigs_T_545; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_547 = _decodeSigs_T_39 ? 4'h0 : _decodeSigs_T_546; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_548 = _decodeSigs_T_37 ? 4'h0 : _decodeSigs_T_547; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_549 = _decodeSigs_T_35 ? 4'h0 : _decodeSigs_T_548; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_550 = _decodeSigs_T_33 ? 4'h0 : _decodeSigs_T_549; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_551 = _decodeSigs_T_31 ? 4'h0 : _decodeSigs_T_550; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_552 = _decodeSigs_T_29 ? 4'h0 : _decodeSigs_T_551; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_553 = _decodeSigs_T_27 ? 4'h0 : _decodeSigs_T_552; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_554 = _decodeSigs_T_25 ? 4'h0 : _decodeSigs_T_553; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_555 = _decodeSigs_T_23 ? 4'h0 : _decodeSigs_T_554; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_556 = _decodeSigs_T_21 ? 4'h0 : _decodeSigs_T_555; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_557 = _decodeSigs_T_19 ? 4'h0 : _decodeSigs_T_556; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_558 = _decodeSigs_T_17 ? 4'h0 : _decodeSigs_T_557; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_559 = _decodeSigs_T_15 ? 4'h0 : _decodeSigs_T_558; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_560 = _decodeSigs_T_13 ? 4'h0 : _decodeSigs_T_559; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_561 = _decodeSigs_T_11 ? 4'h0 : _decodeSigs_T_560; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_562 = _decodeSigs_T_9 ? 4'h0 : _decodeSigs_T_561; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_563 = _decodeSigs_T_7 ? 4'h0 : _decodeSigs_T_562; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_564 = _decodeSigs_T_5 ? 4'h0 : _decodeSigs_T_563; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_565 = _decodeSigs_T_3 ? 4'h0 : _decodeSigs_T_564; // @[Lookup.scala 34:39]
  assign io_out_brType = _decodeSigs_T_1 ? 4'h0 : _decodeSigs_T_142; // @[Lookup.scala 34:39]
  assign io_out_wbType = _decodeSigs_T_1 ? 3'h2 : _decodeSigs_T_189; // @[Lookup.scala 34:39]
  assign io_out_lsuOp = _decodeSigs_T_1 ? 5'h1 : _decodeSigs_T_236; // @[Lookup.scala 34:39]
  assign io_out_aluOp = _decodeSigs_T_1 ? 5'h11 : _decodeSigs_T_283; // @[Lookup.scala 34:39]
  assign io_out_opr1 = _decodeSigs_T_1 ? 4'h1 : _decodeSigs_T_330; // @[Lookup.scala 34:39]
  assign io_out_opr2 = _decodeSigs_T_1 ? 4'h0 : _decodeSigs_T_377; // @[Lookup.scala 34:39]
  assign io_out_immSrc = _decodeSigs_T_1 ? 3'h0 : _decodeSigs_T_424; // @[Lookup.scala 34:39]
  assign io_out_immSign = _decodeSigs_T_1 | (_decodeSigs_T_3 | (_decodeSigs_T_5 | (_decodeSigs_T_7 | (_decodeSigs_T_9 |
    (_decodeSigs_T_11 | _decodeSigs_T_466))))); // @[Lookup.scala 34:39]
  assign io_out_csrOp = _decodeSigs_T_1 ? 3'h0 : _decodeSigs_T_518; // @[Lookup.scala 34:39]
  assign io_out_excpType = _decodeSigs_T_1 ? 4'h0 : _decodeSigs_T_565; // @[Lookup.scala 34:39]
endmodule
module LoadPipe(
  input         clock,
  input         reset,
  output        io_load_req_ready,
  input         io_load_req_valid,
  input  [31:0] io_load_req_bits_addr,
  input         io_load_resp_ready,
  output        io_load_resp_valid,
  output [31:0] io_load_resp_bits_data,
  input         io_dir_req_ready,
  output        io_dir_req_valid,
  output [31:0] io_dir_req_bits_addr,
  input         io_dir_resp_bits_hit,
  input  [3:0]  io_dir_resp_bits_chosenWay,
  input         io_dir_resp_bits_isDirtyWay,
  input  [18:0] io_dir_resp_bits_tagRdVec_0,
  input  [18:0] io_dir_resp_bits_tagRdVec_1,
  input  [18:0] io_dir_resp_bits_tagRdVec_2,
  input  [18:0] io_dir_resp_bits_tagRdVec_3,
  input         io_dataBank_req_ready,
  output        io_dataBank_req_valid,
  output [8:0]  io_dataBank_req_bits_set,
  input  [31:0] io_dataBank_resp_0_0,
  input  [31:0] io_dataBank_resp_0_1,
  input  [31:0] io_dataBank_resp_0_2,
  input  [31:0] io_dataBank_resp_0_3,
  input  [31:0] io_dataBank_resp_1_0,
  input  [31:0] io_dataBank_resp_1_1,
  input  [31:0] io_dataBank_resp_1_2,
  input  [31:0] io_dataBank_resp_1_3,
  input  [31:0] io_dataBank_resp_2_0,
  input  [31:0] io_dataBank_resp_2_1,
  input  [31:0] io_dataBank_resp_2_2,
  input  [31:0] io_dataBank_resp_2_3,
  input  [31:0] io_dataBank_resp_3_0,
  input  [31:0] io_dataBank_resp_3_1,
  input  [31:0] io_dataBank_resp_3_2,
  input  [31:0] io_dataBank_resp_3_3,
  input         io_mshr_ready,
  output        io_mshr_valid,
  output [31:0] io_mshr_bits_addr,
  output        io_mshr_bits_dirInfo_hit,
  output [3:0]  io_mshr_bits_dirInfo_chosenWay,
  output        io_mshr_bits_dirInfo_isDirtyWay,
  output [18:0] io_mshr_bits_dirtyTag,
  output [31:0] io_mshr_bits_data_0,
  output [31:0] io_mshr_bits_data_1,
  output [31:0] io_mshr_bits_data_2,
  output [31:0] io_mshr_bits_data_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  reg  s0_full; // @[LoadPipe.scala 31:26]
  wire  s0_latch = io_load_req_ready & io_load_req_valid; // @[Decoupled.scala 51:35]
  reg  s0_valid_REG; // @[LoadPipe.scala 55:25]
  reg  s0_validReg; // @[LoadPipe.scala 52:30]
  wire  _s0_valid_T_1 = io_dir_req_ready & io_dir_req_valid; // @[Decoupled.scala 51:35]
  wire  _s0_valid_T_3 = io_dataBank_req_ready & io_dataBank_req_valid; // @[Decoupled.scala 51:35]
  wire  s0_valid = (s0_valid_REG | s0_validReg) & _s0_valid_T_1 & _s0_valid_T_3; // @[LoadPipe.scala 55:71]
  reg  s1_full; // @[LoadPipe.scala 61:26]
  reg  s1_dirInfo_hit; // @[Reg.scala 19:16]
  wire  _s1_valid_T = ~s1_dirInfo_hit; // @[LoadPipe.scala 92:21]
  wire  _s1_valid_T_1 = io_mshr_ready & io_mshr_valid; // @[Decoupled.scala 51:35]
  wire  _s1_valid_T_3 = io_load_resp_ready & io_load_resp_valid; // @[Decoupled.scala 51:35]
  wire  _s1_valid_T_4 = s1_dirInfo_hit & _s1_valid_T_3; // @[LoadPipe.scala 93:30]
  wire  _s1_valid_T_5 = ~s1_dirInfo_hit & _s1_valid_T_1 | _s1_valid_T_4; // @[LoadPipe.scala 92:47]
  wire  s1_fire = s1_full & _s1_valid_T_5; // @[LoadPipe.scala 91:25]
  wire  s1_ready = ~s1_full | s1_fire; // @[LoadPipe.scala 75:26]
  wire  s0_fire = s0_valid & s1_ready; // @[LoadPipe.scala 33:28]
  reg [31:0] s0_reqReg_addr; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = s0_latch ? io_load_req_bits_addr : s0_reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_1 = s0_full & s0_fire ? 1'h0 : s0_full; // @[LoadPipe.scala 31:26 40:{35,45}]
  wire  _GEN_2 = s0_latch | _GEN_1; // @[LoadPipe.scala 39:{20,30}]
  wire  _GEN_3 = s0_fire ? 1'h0 : s0_validReg; // @[LoadPipe.scala 54:24 52:30 54:38]
  wire  _GEN_4 = s0_latch | _GEN_3; // @[LoadPipe.scala 53:{20,34}]
  reg [31:0] s1_rAddr; // @[Reg.scala 19:16]
  wire [3:0] s1_blockSel = 4'h1 << s1_rAddr[3:2]; // @[OneHot.scala 57:35]
  reg [31:0] s1_rdDataAll_0_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_3; // @[Reg.scala 19:16]
  reg [3:0] s1_dirInfo_chosenWay; // @[Reg.scala 19:16]
  reg  s1_dirInfo_isDirtyWay; // @[Reg.scala 19:16]
  wire [31:0] _s1_rdBlockData_T_4 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_5 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_6 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_7 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_8 = _s1_rdBlockData_T_4 | _s1_rdBlockData_T_5; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_9 = _s1_rdBlockData_T_8 | _s1_rdBlockData_T_6; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_0 = _s1_rdBlockData_T_9 | _s1_rdBlockData_T_7; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_11 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_12 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_13 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_14 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_15 = _s1_rdBlockData_T_11 | _s1_rdBlockData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_16 = _s1_rdBlockData_T_15 | _s1_rdBlockData_T_13; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_1 = _s1_rdBlockData_T_16 | _s1_rdBlockData_T_14; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_18 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_19 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_20 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_21 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_22 = _s1_rdBlockData_T_18 | _s1_rdBlockData_T_19; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_23 = _s1_rdBlockData_T_22 | _s1_rdBlockData_T_20; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_2 = _s1_rdBlockData_T_23 | _s1_rdBlockData_T_21; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_25 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_26 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_27 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_28 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_29 = _s1_rdBlockData_T_25 | _s1_rdBlockData_T_26; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_30 = _s1_rdBlockData_T_29 | _s1_rdBlockData_T_27; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_3 = _s1_rdBlockData_T_30 | _s1_rdBlockData_T_28; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_4 = s1_blockSel[0] ? s1_rdBlockData_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_5 = s1_blockSel[1] ? s1_rdBlockData_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_6 = s1_blockSel[2] ? s1_rdBlockData_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_7 = s1_blockSel[3] ? s1_rdBlockData_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_8 = _s1_rdData_T_4 | _s1_rdData_T_5; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_9 = _s1_rdData_T_8 | _s1_rdData_T_6; // @[Mux.scala 27:73]
  reg [18:0] s1_tagRdVec_0; // @[Reg.scala 19:16]
  reg [18:0] s1_tagRdVec_1; // @[Reg.scala 19:16]
  reg [18:0] s1_tagRdVec_2; // @[Reg.scala 19:16]
  reg [18:0] s1_tagRdVec_3; // @[Reg.scala 19:16]
  wire [18:0] _s1_dirtyTag_T_4 = s1_dirInfo_chosenWay[0] ? s1_tagRdVec_0 : 19'h0; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_5 = s1_dirInfo_chosenWay[1] ? s1_tagRdVec_1 : 19'h0; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_6 = s1_dirInfo_chosenWay[2] ? s1_tagRdVec_2 : 19'h0; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_7 = s1_dirInfo_chosenWay[3] ? s1_tagRdVec_3 : 19'h0; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_8 = _s1_dirtyTag_T_4 | _s1_dirtyTag_T_5; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_9 = _s1_dirtyTag_T_8 | _s1_dirtyTag_T_6; // @[Mux.scala 27:73]
  wire  _GEN_33 = s1_full & s1_fire ? 1'h0 : s1_full; // @[LoadPipe.scala 61:26 77:{35,45}]
  wire  _GEN_34 = s0_fire | _GEN_33; // @[LoadPipe.scala 76:{20,30}]
  assign io_load_req_ready = ~s0_full; // @[LoadPipe.scala 37:26]
  assign io_load_resp_valid = s1_dirInfo_hit & s1_full; // @[LoadPipe.scala 87:36]
  assign io_load_resp_bits_data = _s1_rdData_T_9 | _s1_rdData_T_7; // @[Mux.scala 27:73]
  assign io_dir_req_valid = s0_latch | s0_full; // @[LoadPipe.scala 43:34]
  assign io_dir_req_bits_addr = s0_latch ? io_load_req_bits_addr : s0_reqReg_addr; // @[LoadPipe.scala 35:23]
  assign io_dataBank_req_valid = s0_latch | s0_full; // @[LoadPipe.scala 46:39]
  assign io_dataBank_req_bits_set = _GEN_0[12:4]; // @[Parameters.scala 50:11]
  assign io_mshr_valid = _s1_valid_T & s1_full; // @[LoadPipe.scala 79:32]
  assign io_mshr_bits_addr = s1_rAddr; // @[LoadPipe.scala 81:23]
  assign io_mshr_bits_dirInfo_hit = s1_dirInfo_hit; // @[LoadPipe.scala 84:26]
  assign io_mshr_bits_dirInfo_chosenWay = s1_dirInfo_chosenWay; // @[LoadPipe.scala 84:26]
  assign io_mshr_bits_dirInfo_isDirtyWay = s1_dirInfo_isDirtyWay; // @[LoadPipe.scala 84:26]
  assign io_mshr_bits_dirtyTag = _s1_dirtyTag_T_9 | _s1_dirtyTag_T_7; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_0 = _s1_rdBlockData_T_9 | _s1_rdBlockData_T_7; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_1 = _s1_rdBlockData_T_16 | _s1_rdBlockData_T_14; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_2 = _s1_rdBlockData_T_23 | _s1_rdBlockData_T_21; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_3 = _s1_rdBlockData_T_30 | _s1_rdBlockData_T_28; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[LoadPipe.scala 31:26]
      s0_full <= 1'h0; // @[LoadPipe.scala 31:26]
    end else begin
      s0_full <= _GEN_2;
    end
    s0_valid_REG <= io_load_req_ready & io_load_req_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[LoadPipe.scala 52:30]
      s0_validReg <= 1'h0; // @[LoadPipe.scala 52:30]
    end else begin
      s0_validReg <= _GEN_4;
    end
    if (reset) begin // @[LoadPipe.scala 61:26]
      s1_full <= 1'h0; // @[LoadPipe.scala 61:26]
    end else begin
      s1_full <= _GEN_34;
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_hit <= io_dir_resp_bits_hit; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_addr <= io_load_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      if (s0_latch) begin // @[Reg.scala 20:18]
        s1_rAddr <= io_load_req_bits_addr; // @[Reg.scala 20:22]
      end else begin
        s1_rAddr <= s0_reqReg_addr; // @[Reg.scala 19:16]
      end
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_0 <= io_dataBank_resp_0_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_1 <= io_dataBank_resp_0_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_2 <= io_dataBank_resp_0_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_3 <= io_dataBank_resp_0_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_0 <= io_dataBank_resp_1_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_1 <= io_dataBank_resp_1_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_2 <= io_dataBank_resp_1_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_3 <= io_dataBank_resp_1_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_0 <= io_dataBank_resp_2_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_1 <= io_dataBank_resp_2_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_2 <= io_dataBank_resp_2_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_3 <= io_dataBank_resp_2_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_0 <= io_dataBank_resp_3_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_1 <= io_dataBank_resp_3_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_2 <= io_dataBank_resp_3_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_3 <= io_dataBank_resp_3_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_chosenWay <= io_dir_resp_bits_chosenWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_isDirtyWay <= io_dir_resp_bits_isDirtyWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_0 <= io_dir_resp_bits_tagRdVec_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_1 <= io_dir_resp_bits_tagRdVec_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_2 <= io_dir_resp_bits_tagRdVec_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_3 <= io_dir_resp_bits_tagRdVec_3; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s0_valid_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s0_validReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s1_full = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s1_dirInfo_hit = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s0_reqReg_addr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  s1_rAddr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  s1_rdDataAll_0_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  s1_rdDataAll_0_1 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  s1_rdDataAll_0_2 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  s1_rdDataAll_0_3 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  s1_rdDataAll_1_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  s1_rdDataAll_1_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  s1_rdDataAll_1_2 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  s1_rdDataAll_1_3 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  s1_rdDataAll_2_0 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  s1_rdDataAll_2_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  s1_rdDataAll_2_2 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  s1_rdDataAll_2_3 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  s1_rdDataAll_3_0 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  s1_rdDataAll_3_1 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  s1_rdDataAll_3_2 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  s1_rdDataAll_3_3 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  s1_dirInfo_chosenWay = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  s1_dirInfo_isDirtyWay = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  s1_tagRdVec_0 = _RAND_25[18:0];
  _RAND_26 = {1{`RANDOM}};
  s1_tagRdVec_1 = _RAND_26[18:0];
  _RAND_27 = {1{`RANDOM}};
  s1_tagRdVec_2 = _RAND_27[18:0];
  _RAND_28 = {1{`RANDOM}};
  s1_tagRdVec_3 = _RAND_28[18:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StorePipe(
  input         clock,
  input         reset,
  output        io_store_req_ready,
  input         io_store_req_valid,
  input  [31:0] io_store_req_bits_addr,
  input  [31:0] io_store_req_bits_data,
  input  [3:0]  io_store_req_bits_mask,
  input         io_store_resp_ready,
  output        io_store_resp_valid,
  output        io_dir_read_req_valid,
  output [31:0] io_dir_read_req_bits_addr,
  input         io_dir_read_resp_bits_hit,
  input  [3:0]  io_dir_read_resp_bits_chosenWay,
  input         io_dir_read_resp_bits_isDirtyWay,
  input  [18:0] io_dir_read_resp_bits_tagRdVec_0,
  input  [18:0] io_dir_read_resp_bits_tagRdVec_1,
  input  [18:0] io_dir_read_resp_bits_tagRdVec_2,
  input  [18:0] io_dir_read_resp_bits_tagRdVec_3,
  output        io_dir_write_req_valid,
  output [31:0] io_dir_write_req_bits_addr,
  output [3:0]  io_dir_write_req_bits_way,
  output        io_dataBank_read_req_valid,
  output [8:0]  io_dataBank_read_req_bits_set,
  input  [31:0] io_dataBank_read_resp_0_0,
  input  [31:0] io_dataBank_read_resp_0_1,
  input  [31:0] io_dataBank_read_resp_0_2,
  input  [31:0] io_dataBank_read_resp_0_3,
  input  [31:0] io_dataBank_read_resp_1_0,
  input  [31:0] io_dataBank_read_resp_1_1,
  input  [31:0] io_dataBank_read_resp_1_2,
  input  [31:0] io_dataBank_read_resp_1_3,
  input  [31:0] io_dataBank_read_resp_2_0,
  input  [31:0] io_dataBank_read_resp_2_1,
  input  [31:0] io_dataBank_read_resp_2_2,
  input  [31:0] io_dataBank_read_resp_2_3,
  input  [31:0] io_dataBank_read_resp_3_0,
  input  [31:0] io_dataBank_read_resp_3_1,
  input  [31:0] io_dataBank_read_resp_3_2,
  input  [31:0] io_dataBank_read_resp_3_3,
  output        io_dataBank_write_req_valid,
  output [8:0]  io_dataBank_write_req_bits_set,
  output [31:0] io_dataBank_write_req_bits_data_0,
  output [31:0] io_dataBank_write_req_bits_data_1,
  output [31:0] io_dataBank_write_req_bits_data_2,
  output [31:0] io_dataBank_write_req_bits_data_3,
  output [3:0]  io_dataBank_write_req_bits_blockMask,
  output [3:0]  io_dataBank_write_req_bits_way,
  input         io_mshr_ready,
  output        io_mshr_valid,
  output [31:0] io_mshr_bits_addr,
  output        io_mshr_bits_dirInfo_hit,
  output [3:0]  io_mshr_bits_dirInfo_chosenWay,
  output        io_mshr_bits_dirInfo_isDirtyWay,
  output [18:0] io_mshr_bits_dirtyTag,
  output [31:0] io_mshr_bits_data_0,
  output [31:0] io_mshr_bits_data_1,
  output [31:0] io_mshr_bits_data_2,
  output [31:0] io_mshr_bits_data_3,
  output [31:0] io_mshr_bits_storeData,
  output [3:0]  io_mshr_bits_storeMask,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  reg  s0_full; // @[StorePipe.scala 31:26]
  wire  s0_latch = io_store_req_ready & io_store_req_valid; // @[Decoupled.scala 51:35]
  reg  s0_valid_REG; // @[StorePipe.scala 57:25]
  reg  s0_validReg; // @[StorePipe.scala 54:30]
  wire  s0_valid = (s0_valid_REG | s0_validReg) & io_dir_read_req_valid & io_dataBank_read_req_valid; // @[StorePipe.scala 57:77]
  reg  s1_full; // @[StorePipe.scala 64:26]
  reg  s1_dirInfo_hit; // @[Reg.scala 19:16]
  wire  _s1_valid_T = ~s1_dirInfo_hit; // @[StorePipe.scala 115:21]
  wire  _s1_valid_T_1 = io_mshr_ready & io_mshr_valid; // @[Decoupled.scala 51:35]
  wire  _s1_valid_T_6 = s1_dirInfo_hit & io_dataBank_write_req_valid & io_dir_write_req_valid; // @[StorePipe.scala 116:60]
  wire  _s1_valid_T_7 = ~s1_dirInfo_hit & _s1_valid_T_1 | _s1_valid_T_6; // @[StorePipe.scala 115:47]
  wire  s1_valid = s1_full & _s1_valid_T_7; // @[StorePipe.scala 114:25]
  reg  s2_full; // @[StorePipe.scala 122:26]
  wire  _s2_valid_T = io_store_resp_ready & io_store_resp_valid; // @[Decoupled.scala 51:35]
  reg  s2_isHit; // @[Reg.scala 19:16]
  wire  s2_fire = _s2_valid_T & s2_full & s2_isHit | ~s2_isHit; // @[StorePipe.scala 134:59]
  wire  s2_ready = ~s2_full | s2_fire; // @[StorePipe.scala 127:26]
  wire  s1_fire = s1_valid & s2_ready; // @[StorePipe.scala 66:28]
  wire  s1_ready = (~s1_full | s1_fire) & io_mshr_ready; // @[StorePipe.scala 81:39]
  wire  s0_fire = s0_valid & s1_ready; // @[StorePipe.scala 33:28]
  reg [31:0] s0_reqReg_addr; // @[Reg.scala 19:16]
  reg [31:0] s0_reqReg_data; // @[Reg.scala 19:16]
  reg [3:0] s0_reqReg_mask; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = s0_latch ? io_store_req_bits_addr : s0_reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_3 = s0_full & s0_fire ? 1'h0 : s0_full; // @[StorePipe.scala 31:26 41:{35,45}]
  wire  _GEN_4 = s0_latch | _GEN_3; // @[StorePipe.scala 40:{20,30}]
  wire  _GEN_5 = s0_fire ? 1'h0 : s0_validReg; // @[StorePipe.scala 56:24 54:30 56:38]
  wire  _GEN_6 = s0_latch | _GEN_5; // @[StorePipe.scala 55:{20,34}]
  reg [31:0] s1_reqReg_addr; // @[Reg.scala 19:16]
  reg [31:0] s1_reqReg_data; // @[Reg.scala 19:16]
  reg [3:0] s1_reqReg_mask; // @[Reg.scala 19:16]
  wire [3:0] s1_dataBlockSelOH = 4'h1 << s1_reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  reg [31:0] s1_rdDataAll_0_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_3; // @[Reg.scala 19:16]
  reg [3:0] s1_dirInfo_chosenWay; // @[Reg.scala 19:16]
  reg  s1_dirInfo_isDirtyWay; // @[Reg.scala 19:16]
  wire [31:0] _s1_rdBlockData_T_4 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_5 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_6 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_7 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_8 = _s1_rdBlockData_T_4 | _s1_rdBlockData_T_5; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_9 = _s1_rdBlockData_T_8 | _s1_rdBlockData_T_6; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_0 = _s1_rdBlockData_T_9 | _s1_rdBlockData_T_7; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_11 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_12 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_13 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_14 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_15 = _s1_rdBlockData_T_11 | _s1_rdBlockData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_16 = _s1_rdBlockData_T_15 | _s1_rdBlockData_T_13; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_1 = _s1_rdBlockData_T_16 | _s1_rdBlockData_T_14; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_18 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_19 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_20 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_21 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_22 = _s1_rdBlockData_T_18 | _s1_rdBlockData_T_19; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_23 = _s1_rdBlockData_T_22 | _s1_rdBlockData_T_20; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_2 = _s1_rdBlockData_T_23 | _s1_rdBlockData_T_21; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_25 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_26 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_27 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_28 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_29 = _s1_rdBlockData_T_25 | _s1_rdBlockData_T_26; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_30 = _s1_rdBlockData_T_29 | _s1_rdBlockData_T_27; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_3 = _s1_rdBlockData_T_30 | _s1_rdBlockData_T_28; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_4 = s1_dataBlockSelOH[0] ? s1_rdBlockData_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_5 = s1_dataBlockSelOH[1] ? s1_rdBlockData_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_6 = s1_dataBlockSelOH[2] ? s1_rdBlockData_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_7 = s1_dataBlockSelOH[3] ? s1_rdBlockData_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_8 = _s1_rdData_T_4 | _s1_rdData_T_5; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_9 = _s1_rdData_T_8 | _s1_rdData_T_6; // @[Mux.scala 27:73]
  wire [31:0] s1_rdData = _s1_rdData_T_9 | _s1_rdData_T_7; // @[Mux.scala 27:73]
  reg [18:0] s1_tagRdVec_0; // @[Reg.scala 19:16]
  reg [18:0] s1_tagRdVec_1; // @[Reg.scala 19:16]
  reg [18:0] s1_tagRdVec_2; // @[Reg.scala 19:16]
  reg [18:0] s1_tagRdVec_3; // @[Reg.scala 19:16]
  wire [18:0] _s1_dirtyTag_T_4 = s1_dirInfo_chosenWay[0] ? s1_tagRdVec_0 : 19'h0; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_5 = s1_dirInfo_chosenWay[1] ? s1_tagRdVec_1 : 19'h0; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_6 = s1_dirInfo_chosenWay[2] ? s1_tagRdVec_2 : 19'h0; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_7 = s1_dirInfo_chosenWay[3] ? s1_tagRdVec_3 : 19'h0; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_8 = _s1_dirtyTag_T_4 | _s1_dirtyTag_T_5; // @[Mux.scala 27:73]
  wire [18:0] _s1_dirtyTag_T_9 = _s1_dirtyTag_T_8 | _s1_dirtyTag_T_6; // @[Mux.scala 27:73]
  wire  _GEN_37 = s1_full & s1_fire ? 1'h0 : s1_full; // @[StorePipe.scala 64:26 83:{35,45}]
  wire  _GEN_38 = s0_fire | _GEN_37; // @[StorePipe.scala 82:{20,30}]
  wire [1:0] hi = s1_dataBlockSelOH[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo = s1_dataBlockSelOH[1:0]; // @[OneHot.scala 31:18]
  wire  _T_2 = |hi; // @[OneHot.scala 32:14]
  wire [1:0] _T_3 = hi | lo; // @[OneHot.scala 32:28]
  wire [1:0] _T_5 = {_T_2,_T_3[1]}; // @[Cat.scala 33:92]
  wire [7:0] _tempWrData_tempMask_T_5 = s1_reqReg_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_7 = s1_reqReg_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_9 = s1_reqReg_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_11 = s1_reqReg_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [31:0] tempWrData_tempMask = {_tempWrData_tempMask_T_11,_tempWrData_tempMask_T_9,_tempWrData_tempMask_T_7,
    _tempWrData_tempMask_T_5}; // @[Cat.scala 33:92]
  wire [31:0] _tempWrData_T = ~tempWrData_tempMask; // @[Parameters.scala 67:8]
  wire [31:0] _tempWrData_T_1 = _tempWrData_T & s1_rdData; // @[Parameters.scala 67:18]
  wire [31:0] _tempWrData_T_2 = tempWrData_tempMask & s1_reqReg_data; // @[Parameters.scala 67:41]
  wire [31:0] _tempWrData_T_3 = _tempWrData_T_1 | _tempWrData_T_2; // @[Parameters.scala 67:29]
  wire  _GEN_44 = s2_full & s2_fire ? 1'h0 : s2_full; // @[StorePipe.scala 122:26 129:{35,45}]
  wire  _GEN_45 = s1_fire | _GEN_44; // @[StorePipe.scala 128:{20,30}]
  assign io_store_req_ready = ~s0_full; // @[StorePipe.scala 39:27]
  assign io_store_resp_valid = s2_isHit & s2_full & ~io_flush; // @[StorePipe.scala 131:48]
  assign io_dir_read_req_valid = s0_latch | s0_full; // @[StorePipe.scala 44:39]
  assign io_dir_read_req_bits_addr = s0_latch ? io_store_req_bits_addr : s0_reqReg_addr; // @[StorePipe.scala 35:23]
  assign io_dir_write_req_valid = s1_dirInfo_hit & s1_full; // @[StorePipe.scala 95:40]
  assign io_dir_write_req_bits_addr = s1_reqReg_addr; // @[StorePipe.scala 97:32]
  assign io_dir_write_req_bits_way = s1_dirInfo_chosenWay; // @[StorePipe.scala 102:31]
  assign io_dataBank_read_req_valid = s0_latch | s0_full; // @[StorePipe.scala 47:44]
  assign io_dataBank_read_req_bits_set = _GEN_0[12:4]; // @[Parameters.scala 50:11]
  assign io_dataBank_write_req_valid = s1_dirInfo_hit & s1_full; // @[StorePipe.scala 104:45]
  assign io_dataBank_write_req_bits_set = s1_reqReg_addr[12:4]; // @[Parameters.scala 50:11]
  assign io_dataBank_write_req_bits_data_0 = 2'h0 == _T_5 ? _tempWrData_T_3 : 32'h0; // @[StorePipe.scala 109:30 110:{45,45}]
  assign io_dataBank_write_req_bits_data_1 = 2'h1 == _T_5 ? _tempWrData_T_3 : 32'h0; // @[StorePipe.scala 109:30 110:{45,45}]
  assign io_dataBank_write_req_bits_data_2 = 2'h2 == _T_5 ? _tempWrData_T_3 : 32'h0; // @[StorePipe.scala 109:30 110:{45,45}]
  assign io_dataBank_write_req_bits_data_3 = 2'h3 == _T_5 ? _tempWrData_T_3 : 32'h0; // @[StorePipe.scala 109:30 110:{45,45}]
  assign io_dataBank_write_req_bits_blockMask = 4'h1 << s1_reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  assign io_dataBank_write_req_bits_way = s1_dirInfo_chosenWay; // @[StorePipe.scala 108:36]
  assign io_mshr_valid = _s1_valid_T & s1_full; // @[StorePipe.scala 85:32]
  assign io_mshr_bits_addr = s1_reqReg_addr; // @[StorePipe.scala 87:23]
  assign io_mshr_bits_dirInfo_hit = s1_dirInfo_hit; // @[StorePipe.scala 88:26]
  assign io_mshr_bits_dirInfo_chosenWay = s1_dirInfo_chosenWay; // @[StorePipe.scala 88:26]
  assign io_mshr_bits_dirInfo_isDirtyWay = s1_dirInfo_isDirtyWay; // @[StorePipe.scala 88:26]
  assign io_mshr_bits_dirtyTag = _s1_dirtyTag_T_9 | _s1_dirtyTag_T_7; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_0 = _s1_rdBlockData_T_9 | _s1_rdBlockData_T_7; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_1 = _s1_rdBlockData_T_16 | _s1_rdBlockData_T_14; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_2 = _s1_rdBlockData_T_23 | _s1_rdBlockData_T_21; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_3 = _s1_rdBlockData_T_30 | _s1_rdBlockData_T_28; // @[Mux.scala 27:73]
  assign io_mshr_bits_storeData = s1_reqReg_data; // @[StorePipe.scala 92:28]
  assign io_mshr_bits_storeMask = s1_reqReg_mask; // @[StorePipe.scala 93:28]
  always @(posedge clock) begin
    if (reset) begin // @[StorePipe.scala 31:26]
      s0_full <= 1'h0; // @[StorePipe.scala 31:26]
    end else if (io_flush) begin // @[StorePipe.scala 136:20]
      s0_full <= 1'h0; // @[StorePipe.scala 137:17]
    end else begin
      s0_full <= _GEN_4;
    end
    s0_valid_REG <= io_store_req_ready & io_store_req_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[StorePipe.scala 54:30]
      s0_validReg <= 1'h0; // @[StorePipe.scala 54:30]
    end else begin
      s0_validReg <= _GEN_6;
    end
    if (reset) begin // @[StorePipe.scala 64:26]
      s1_full <= 1'h0; // @[StorePipe.scala 64:26]
    end else if (io_flush) begin // @[StorePipe.scala 136:20]
      s1_full <= 1'h0; // @[StorePipe.scala 138:17]
    end else begin
      s1_full <= _GEN_38;
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_hit <= io_dir_read_resp_bits_hit; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[StorePipe.scala 122:26]
      s2_full <= 1'h0; // @[StorePipe.scala 122:26]
    end else if (io_flush) begin // @[StorePipe.scala 136:20]
      s2_full <= 1'h0; // @[StorePipe.scala 139:17]
    end else begin
      s2_full <= _GEN_45;
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_isHit <= s1_dirInfo_hit; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_addr <= io_store_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_data <= io_store_req_bits_data; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_mask <= io_store_req_bits_mask; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_reqReg_addr <= s0_reqReg_addr; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_reqReg_data <= s0_reqReg_data; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_reqReg_mask <= s0_reqReg_mask; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_0 <= io_dataBank_read_resp_0_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_1 <= io_dataBank_read_resp_0_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_2 <= io_dataBank_read_resp_0_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_3 <= io_dataBank_read_resp_0_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_0 <= io_dataBank_read_resp_1_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_1 <= io_dataBank_read_resp_1_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_2 <= io_dataBank_read_resp_1_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_3 <= io_dataBank_read_resp_1_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_0 <= io_dataBank_read_resp_2_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_1 <= io_dataBank_read_resp_2_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_2 <= io_dataBank_read_resp_2_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_3 <= io_dataBank_read_resp_2_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_0 <= io_dataBank_read_resp_3_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_1 <= io_dataBank_read_resp_3_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_2 <= io_dataBank_read_resp_3_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_3 <= io_dataBank_read_resp_3_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_chosenWay <= io_dir_read_resp_bits_chosenWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_isDirtyWay <= io_dir_read_resp_bits_isDirtyWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_0 <= io_dir_read_resp_bits_tagRdVec_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_1 <= io_dir_read_resp_bits_tagRdVec_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_2 <= io_dir_read_resp_bits_tagRdVec_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_3 <= io_dir_read_resp_bits_tagRdVec_3; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s0_valid_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s0_validReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s1_full = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s1_dirInfo_hit = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s2_full = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s2_isHit = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s0_reqReg_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  s0_reqReg_data = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  s0_reqReg_mask = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  s1_reqReg_addr = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  s1_reqReg_data = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  s1_reqReg_mask = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  s1_rdDataAll_0_0 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  s1_rdDataAll_0_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  s1_rdDataAll_0_2 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  s1_rdDataAll_0_3 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  s1_rdDataAll_1_0 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  s1_rdDataAll_1_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  s1_rdDataAll_1_2 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  s1_rdDataAll_1_3 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  s1_rdDataAll_2_0 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  s1_rdDataAll_2_1 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  s1_rdDataAll_2_2 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  s1_rdDataAll_2_3 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  s1_rdDataAll_3_0 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  s1_rdDataAll_3_1 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  s1_rdDataAll_3_2 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  s1_rdDataAll_3_3 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  s1_dirInfo_chosenWay = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  s1_dirInfo_isDirtyWay = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  s1_tagRdVec_0 = _RAND_31[18:0];
  _RAND_32 = {1{`RANDOM}};
  s1_tagRdVec_1 = _RAND_32[18:0];
  _RAND_33 = {1{`RANDOM}};
  s1_tagRdVec_2 = _RAND_33[18:0];
  _RAND_34 = {1{`RANDOM}};
  s1_tagRdVec_3 = _RAND_34[18:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MSHR(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [31:0] io_req_bits_addr,
  input         io_req_bits_dirInfo_hit,
  input  [3:0]  io_req_bits_dirInfo_chosenWay,
  input         io_req_bits_dirInfo_isDirtyWay,
  input  [18:0] io_req_bits_dirtyTag,
  input  [31:0] io_req_bits_data_0,
  input  [31:0] io_req_bits_data_1,
  input  [31:0] io_req_bits_data_2,
  input  [31:0] io_req_bits_data_3,
  input         io_req_bits_isStore,
  input  [31:0] io_req_bits_storeData,
  input  [3:0]  io_req_bits_storeMask,
  input         io_resp_load_ready,
  output        io_resp_load_valid,
  output [31:0] io_resp_load_bits_data,
  input         io_resp_store_ready,
  output        io_resp_store_valid,
  output        io_tasks_refill_req_valid,
  output [31:0] io_tasks_refill_req_bits_addr,
  output [3:0]  io_tasks_refill_req_bits_chosenWay,
  output        io_tasks_refill_resp_ready,
  input         io_tasks_refill_resp_valid,
  input  [31:0] io_tasks_refill_resp_bits_data,
  output        io_tasks_writeback_req_valid,
  output [31:0] io_tasks_writeback_req_bits_addr,
  output [18:0] io_tasks_writeback_req_bits_dirtyTag,
  output [31:0] io_tasks_writeback_req_bits_data_0,
  output [31:0] io_tasks_writeback_req_bits_data_1,
  output [31:0] io_tasks_writeback_req_bits_data_2,
  output [31:0] io_tasks_writeback_req_bits_data_3,
  output        io_tasks_writeback_resp_ready,
  input         io_tasks_writeback_resp_valid,
  input         io_dirWrite_req_ready,
  output        io_dirWrite_req_valid,
  output [31:0] io_dirWrite_req_bits_addr,
  output [3:0]  io_dirWrite_req_bits_way,
  input         io_dataWrite_req_ready,
  output        io_dataWrite_req_valid,
  output [8:0]  io_dataWrite_req_bits_set,
  output [31:0] io_dataWrite_req_bits_data_0,
  output [31:0] io_dataWrite_req_bits_data_1,
  output [31:0] io_dataWrite_req_bits_data_2,
  output [31:0] io_dataWrite_req_bits_data_3,
  output [3:0]  io_dataWrite_req_bits_blockMask,
  output [3:0]  io_dataWrite_req_bits_way,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] reqReg_addr; // @[Reg.scala 19:16]
  reg [3:0] reqReg_dirInfo_chosenWay; // @[Reg.scala 19:16]
  reg [18:0] reqReg_dirtyTag; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_0; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_1; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_2; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_3; // @[Reg.scala 19:16]
  reg  reqReg_isStore; // @[Reg.scala 19:16]
  reg [31:0] reqReg_storeData; // @[Reg.scala 19:16]
  reg [3:0] reqReg_storeMask; // @[Reg.scala 19:16]
  wire  _GEN_13 = _reqReg_T ? io_req_bits_isStore : reqReg_isStore; // @[Reg.scala 19:16 20:{18,22}]
  reg [2:0] state; // @[MSHR.scala 65:24]
  wire  _io_busy_T = state == 3'h0; // @[MSHR.scala 68:22]
  wire [1:0] _GEN_17 = io_req_bits_dirInfo_isDirtyWay ? 2'h1 : 2'h2; // @[MSHR.scala 75:50 76:27 78:27]
  wire [1:0] _GEN_18 = _reqReg_T ? _GEN_17 : 2'h0; // @[MSHR.scala 73:19 74:27]
  wire [1:0] _GEN_19 = _io_busy_T ? _GEN_18 : 2'h0; // @[MSHR.scala 72:27 66:29]
  wire  _T_2 = state == 3'h1; // @[MSHR.scala 84:16]
  wire  _T_3 = io_tasks_writeback_resp_ready & io_tasks_writeback_resp_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_20 = _T_3 ? 2'h2 : 2'h1; // @[MSHR.scala 85:19 86:44 87:23]
  wire [1:0] _GEN_21 = state == 3'h1 ? _GEN_20 : _GEN_19; // @[MSHR.scala 84:32]
  wire  _T_4 = state == 3'h2; // @[MSHR.scala 92:16]
  wire  _T_5 = io_tasks_refill_resp_ready & io_tasks_refill_resp_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_22 = _T_5 ? 3'h4 : 3'h2; // @[MSHR.scala 93:19 96:47 97:23]
  wire [2:0] _GEN_23 = _T_5 & _GEN_13 ? 3'h3 : _GEN_22; // @[MSHR.scala 94:56 95:23]
  wire  _T_8 = io_resp_load_ready & io_resp_load_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_24 = _T_8 ? 3'h0 : _GEN_23; // @[MSHR.scala 100:33 101:23]
  wire [2:0] _GEN_25 = state == 3'h2 ? _GEN_24 : {{1'd0}, _GEN_21}; // @[MSHR.scala 92:29]
  wire  _T_9 = state == 3'h3; // @[MSHR.scala 106:16]
  wire  _T_10 = io_dirWrite_req_ready & io_dirWrite_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_11 = io_dataWrite_req_ready & io_dataWrite_req_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_26 = _T_10 & _T_11 ? 3'h4 : 3'h3; // @[MSHR.scala 107:19 108:61 109:23]
  wire  _T_13 = io_resp_store_ready & io_resp_store_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_27 = _T_13 ? 3'h0 : _GEN_26; // @[MSHR.scala 112:34 113:23]
  wire  _T_14 = state == 3'h4; // @[MSHR.scala 118:16]
  wire  _willRefill_T_1 = ~io_req_bits_dirInfo_hit; // @[MSHR.scala 127:63]
  wire  willRefill = ~io_req_bits_dirInfo_isDirtyWay & ~io_req_bits_dirInfo_hit & _reqReg_T; // @[MSHR.scala 127:88]
  wire  willWriteback = io_req_bits_dirInfo_isDirtyWay & _willRefill_T_1 & _reqReg_T; // @[MSHR.scala 128:87]
  wire  willWriteStore = _T_4 & _GEN_13 & _T_5; // @[MSHR.scala 129:61]
  wire  _willRespLoad_T_1 = ~_GEN_13; // @[MSHR.scala 130:49]
  wire  willRespLoad = _T_4 & ~_GEN_13 & _T_5; // @[MSHR.scala 130:62]
  wire  willRespStore = _T_9 & _T_10 & _T_11; // @[MSHR.scala 131:73]
  wire  _io_dirWrite_req_valid_T_1 = _T_9 | willWriteStore; // @[MSHR.scala 146:51]
  wire  _io_dataWrite_req_valid_T_2 = ~io_flush; // @[MSHR.scala 155:75]
  wire [3:0] _io_dataWrite_req_bits_blockMask_T_1 = 4'h1 << reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  reg [31:0] oldData_r; // @[Reg.scala 19:16]
  wire [31:0] _GEN_31 = _T_5 ? io_tasks_refill_resp_bits_data : oldData_r; // @[Reg.scala 19:16 20:{18,22}]
  wire [1:0] hi = _io_dataWrite_req_bits_blockMask_T_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo = _io_dataWrite_req_bits_blockMask_T_1[1:0]; // @[OneHot.scala 31:18]
  wire  _T_20 = |hi; // @[OneHot.scala 32:14]
  wire [1:0] _T_21 = hi | lo; // @[OneHot.scala 32:28]
  wire [1:0] _T_23 = {_T_20,_T_21[1]}; // @[Cat.scala 33:92]
  wire [7:0] _tempWrData_tempMask_T_5 = reqReg_storeMask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_7 = reqReg_storeMask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_9 = reqReg_storeMask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_11 = reqReg_storeMask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [31:0] tempWrData_tempMask = {_tempWrData_tempMask_T_11,_tempWrData_tempMask_T_9,_tempWrData_tempMask_T_7,
    _tempWrData_tempMask_T_5}; // @[Cat.scala 33:92]
  wire [31:0] _tempWrData_T = ~tempWrData_tempMask; // @[Parameters.scala 67:8]
  wire [31:0] _tempWrData_T_1 = _tempWrData_T & _GEN_31; // @[Parameters.scala 67:18]
  wire [31:0] _tempWrData_T_2 = tempWrData_tempMask & reqReg_storeData; // @[Parameters.scala 67:41]
  wire [31:0] _tempWrData_T_3 = _tempWrData_T_1 | _tempWrData_T_2; // @[Parameters.scala 67:29]
  reg [31:0] io_resp_load_bits_data_r; // @[Reg.scala 19:16]
  assign io_req_ready = state == 3'h0; // @[MSHR.scala 69:27]
  assign io_resp_load_valid = _willRespLoad_T_1 & (_T_14 | willRespLoad) & _io_dataWrite_req_valid_T_2; // @[MSHR.scala 167:77]
  assign io_resp_load_bits_data = _T_5 ? io_tasks_refill_resp_bits_data : io_resp_load_bits_data_r; // @[MSHR.scala 168:34]
  assign io_resp_store_valid = _GEN_13 & (_T_14 | willRespStore); // @[MSHR.scala 173:40]
  assign io_tasks_refill_req_valid = _T_4 | willRefill; // @[MSHR.scala 133:52]
  assign io_tasks_refill_req_bits_addr = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[MSHR.scala 61:18]
  assign io_tasks_refill_req_bits_chosenWay = _reqReg_T ? io_req_bits_dirInfo_chosenWay : reqReg_dirInfo_chosenWay; // @[MSHR.scala 61:18]
  assign io_tasks_refill_resp_ready = 1'h1; // @[MSHR.scala 136:32]
  assign io_tasks_writeback_req_valid = _T_2 | willWriteback; // @[MSHR.scala 139:58]
  assign io_tasks_writeback_req_bits_addr = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[MSHR.scala 61:18]
  assign io_tasks_writeback_req_bits_dirtyTag = _reqReg_T ? io_req_bits_dirtyTag : reqReg_dirtyTag; // @[MSHR.scala 61:18]
  assign io_tasks_writeback_req_bits_data_0 = _reqReg_T ? io_req_bits_data_0 : reqReg_data_0; // @[MSHR.scala 61:18]
  assign io_tasks_writeback_req_bits_data_1 = _reqReg_T ? io_req_bits_data_1 : reqReg_data_1; // @[MSHR.scala 61:18]
  assign io_tasks_writeback_req_bits_data_2 = _reqReg_T ? io_req_bits_data_2 : reqReg_data_2; // @[MSHR.scala 61:18]
  assign io_tasks_writeback_req_bits_data_3 = _reqReg_T ? io_req_bits_data_3 : reqReg_data_3; // @[MSHR.scala 61:18]
  assign io_tasks_writeback_resp_ready = 1'h1; // @[MSHR.scala 143:35]
  assign io_dirWrite_req_valid = _T_9 | willWriteStore; // @[MSHR.scala 146:51]
  assign io_dirWrite_req_bits_addr = reqReg_addr; // @[MSHR.scala 147:31]
  assign io_dirWrite_req_bits_way = reqReg_dirInfo_chosenWay; // @[MSHR.scala 152:30]
  assign io_dataWrite_req_valid = _io_dirWrite_req_valid_T_1 & ~io_flush; // @[MSHR.scala 155:72]
  assign io_dataWrite_req_bits_set = reqReg_addr[12:4]; // @[Parameters.scala 50:11]
  assign io_dataWrite_req_bits_data_0 = 2'h0 == _T_23 ? _tempWrData_T_3 : 32'h0; // @[MSHR.scala 160:30 161:{60,60}]
  assign io_dataWrite_req_bits_data_1 = 2'h1 == _T_23 ? _tempWrData_T_3 : 32'h0; // @[MSHR.scala 160:30 161:{60,60}]
  assign io_dataWrite_req_bits_data_2 = 2'h2 == _T_23 ? _tempWrData_T_3 : 32'h0; // @[MSHR.scala 160:30 161:{60,60}]
  assign io_dataWrite_req_bits_data_3 = 2'h3 == _T_23 ? _tempWrData_T_3 : 32'h0; // @[MSHR.scala 160:30 161:{60,60}]
  assign io_dataWrite_req_bits_blockMask = 4'h1 << reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  assign io_dataWrite_req_bits_way = reqReg_dirInfo_chosenWay; // @[MSHR.scala 158:31]
  always @(posedge clock) begin
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_addr <= io_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_dirInfo_chosenWay <= io_req_bits_dirInfo_chosenWay; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_dirtyTag <= io_req_bits_dirtyTag; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_0 <= io_req_bits_data_0; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_1 <= io_req_bits_data_1; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_2 <= io_req_bits_data_2; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_3 <= io_req_bits_data_3; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_isStore <= io_req_bits_isStore; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_storeData <= io_req_bits_storeData; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_storeMask <= io_req_bits_storeMask; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[MSHR.scala 65:24]
      state <= 3'h0; // @[MSHR.scala 65:24]
    end else if (io_flush) begin // @[MSHR.scala 175:20]
      state <= 3'h0; // @[MSHR.scala 176:15]
    end else if (state == 3'h4) begin // @[MSHR.scala 118:27]
      if (_T_8 | _T_13) begin // @[MSHR.scala 120:55]
        state <= 3'h0; // @[MSHR.scala 121:23]
      end else begin
        state <= 3'h4; // @[MSHR.scala 119:19]
      end
    end else if (state == 3'h3) begin // @[MSHR.scala 106:32]
      state <= _GEN_27;
    end else begin
      state <= _GEN_25;
    end
    if (_T_5) begin // @[Reg.scala 20:18]
      oldData_r <= io_tasks_refill_resp_bits_data; // @[Reg.scala 20:22]
    end
    if (_T_5) begin // @[Reg.scala 20:18]
      io_resp_load_bits_data_r <= io_tasks_refill_resp_bits_data; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reqReg_addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reqReg_dirInfo_chosenWay = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  reqReg_dirtyTag = _RAND_2[18:0];
  _RAND_3 = {1{`RANDOM}};
  reqReg_data_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reqReg_data_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reqReg_data_2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reqReg_data_3 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reqReg_isStore = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reqReg_storeData = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reqReg_storeMask = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  oldData_r = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  io_resp_load_bits_data_r = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RefillPipe_1(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [31:0]  io_req_bits_addr,
  input  [3:0]   io_req_bits_chosenWay,
  output         io_resp_valid,
  output [31:0]  io_resp_bits_data,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [31:0]  io_tlbus_req_bits_address,
  output         io_tlbus_resp_ready,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data,
  input          io_dirWrite_req_ready,
  output         io_dirWrite_req_valid,
  output [31:0]  io_dirWrite_req_bits_addr,
  output [3:0]   io_dirWrite_req_bits_way,
  input          io_dataWrite_req_ready,
  output         io_dataWrite_req_valid,
  output [8:0]   io_dataWrite_req_bits_set,
  output [31:0]  io_dataWrite_req_bits_data_0,
  output [31:0]  io_dataWrite_req_bits_data_1,
  output [31:0]  io_dataWrite_req_bits_data_2,
  output [31:0]  io_dataWrite_req_bits_data_3,
  output [3:0]   io_dataWrite_req_bits_way
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[RefillPipe.scala 42:24]
  wire  _io_req_ready_T = state == 2'h0; // @[RefillPipe.scala 45:27]
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] reqReg_addr; // @[Reg.scala 19:16]
  reg [3:0] reqReg_chosenWay; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  reg  reqValidReg; // @[Reg.scala 19:16]
  wire  _GEN_2 = _reqReg_T | reqValidReg; // @[Reg.scala 19:16 20:{18,22}]
  wire [3:0] dataBlockSelOH = 4'h1 << reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  wire  _refillFire_T = io_tlbus_resp_ready & io_tlbus_resp_valid; // @[Decoupled.scala 51:35]
  wire  refillFire = _refillFire_T & io_tlbus_resp_bits_opcode == 3'h1; // @[RefillPipe.scala 59:41]
  wire  _T_2 = io_tlbus_req_ready & io_tlbus_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_4 = _T_2 ? 2'h2 : {{1'd0}, _reqReg_T}; // @[RefillPipe.scala 71:33 72:23]
  wire  _GEN_5 = _T_2 ? 1'h0 : _GEN_2; // @[RefillPipe.scala 71:33 73:25]
  wire [1:0] _GEN_6 = _io_req_ready_T ? _GEN_4 : 2'h0; // @[RefillPipe.scala 66:27 43:29]
  wire  _GEN_7 = _io_req_ready_T ? _GEN_5 : _GEN_2; // @[RefillPipe.scala 66:27]
  wire [1:0] _GEN_8 = _T_2 ? 2'h2 : 2'h1; // @[RefillPipe.scala 80:19 81:33 82:23]
  wire  _T_5 = state == 2'h2; // @[RefillPipe.scala 89:16]
  wire [1:0] _GEN_12 = io_resp_valid ? 2'h0 : 2'h3; // @[RefillPipe.scala 92:23 93:32 94:27]
  wire  _T_7 = state == 2'h3; // @[RefillPipe.scala 105:16]
  wire [31:0] _io_resp_bits_data_T_8 = dataBlockSelOH[0] ? io_tlbus_resp_bits_data[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_9 = dataBlockSelOH[1] ? io_tlbus_resp_bits_data[63:32] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_10 = dataBlockSelOH[2] ? io_tlbus_resp_bits_data[95:64] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_11 = dataBlockSelOH[3] ? io_tlbus_resp_bits_data[127:96] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_12 = _io_resp_bits_data_T_8 | _io_resp_bits_data_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_13 = _io_resp_bits_data_T_12 | _io_resp_bits_data_T_10; // @[Mux.scala 27:73]
  assign io_req_ready = state == 2'h0; // @[RefillPipe.scala 45:27]
  assign io_resp_valid = _T_7 | refillFire; // @[RefillPipe.scala 140:38]
  assign io_resp_bits_data = _io_resp_bits_data_T_13 | _io_resp_bits_data_T_11; // @[Mux.scala 27:73]
  assign io_tlbus_req_valid = _reqReg_T | reqValidReg; // @[RefillPipe.scala 50:23]
  assign io_tlbus_req_bits_address = {_GEN_0[31:4],4'h0}; // @[Cat.scala 33:92]
  assign io_tlbus_resp_ready = io_dataWrite_req_ready & io_dirWrite_req_ready; // @[RefillPipe.scala 62:51]
  assign io_dirWrite_req_valid = refillFire & _T_5; // @[RefillPipe.scala 115:33]
  assign io_dirWrite_req_bits_addr = reqReg_addr; // @[RefillPipe.scala 117:31]
  assign io_dirWrite_req_bits_way = reqReg_chosenWay; // @[RefillPipe.scala 122:30]
  assign io_dataWrite_req_valid = refillFire & _T_5; // @[RefillPipe.scala 115:33]
  assign io_dataWrite_req_bits_set = reqReg_addr[12:4]; // @[Parameters.scala 50:11]
  assign io_dataWrite_req_bits_data_0 = io_tlbus_resp_bits_data[31:0]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_1 = io_tlbus_resp_bits_data[63:32]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_2 = io_tlbus_resp_bits_data[95:64]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_3 = io_tlbus_resp_bits_data[127:96]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_way = reqReg_chosenWay; // @[RefillPipe.scala 128:31]
  always @(posedge clock) begin
    if (reset) begin // @[RefillPipe.scala 42:24]
      state <= 2'h0; // @[RefillPipe.scala 42:24]
    end else if (state == 2'h3) begin // @[RefillPipe.scala 105:27]
      state <= _GEN_12;
    end else if (state == 2'h2) begin // @[RefillPipe.scala 89:33]
      if (refillFire) begin // @[RefillPipe.scala 91:30]
        state <= _GEN_12;
      end else begin
        state <= 2'h2;
      end
    end else if (state == 2'h1) begin // @[RefillPipe.scala 79:26]
      state <= _GEN_8;
    end else begin
      state <= _GEN_6;
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_addr <= io_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_chosenWay <= io_req_bits_chosenWay; // @[Reg.scala 20:22]
    end
    if (state == 2'h1) begin // @[RefillPipe.scala 79:26]
      if (_T_2) begin // @[RefillPipe.scala 81:33]
        reqValidReg <= 1'h0; // @[RefillPipe.scala 83:25]
      end else begin
        reqValidReg <= _GEN_7;
      end
    end else begin
      reqValidReg <= _GEN_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reqReg_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqReg_chosenWay = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  reqValidReg = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLSerializer(
  input         io_in_valid,
  input  [31:0] io_in_bits_0_0,
  input  [31:0] io_in_bits_0_1,
  input  [31:0] io_in_bits_0_2,
  input  [31:0] io_in_bits_0_3,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_0,
  output [31:0] io_out_bits_1,
  output [31:0] io_out_bits_2,
  output [31:0] io_out_bits_3,
  output        io_fireAll
);
  assign io_out_valid = io_in_valid; // @[TLSerializer.scala 41:18]
  assign io_out_bits_0 = io_in_bits_0_0; // @[TLSerializer.scala 42:17]
  assign io_out_bits_1 = io_in_bits_0_1; // @[TLSerializer.scala 42:17]
  assign io_out_bits_2 = io_in_bits_0_2; // @[TLSerializer.scala 42:17]
  assign io_out_bits_3 = io_in_bits_0_3; // @[TLSerializer.scala 42:17]
  assign io_fireAll = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
endmodule
module WritebackQueue(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [31:0]  io_req_bits_addr,
  input  [18:0]  io_req_bits_dirtyTag,
  input  [31:0]  io_req_bits_data_0,
  input  [31:0]  io_req_bits_data_1,
  input  [31:0]  io_req_bits_data_2,
  input  [31:0]  io_req_bits_data_3,
  output         io_resp_valid,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [31:0]  io_tlbus_req_bits_address,
  output [127:0] io_tlbus_req_bits_data,
  output         io_tlbus_resp_ready,
  input          io_tlbus_resp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  serializer_io_in_valid; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_in_bits_0_0; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_in_bits_0_1; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_in_bits_0_2; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_in_bits_0_3; // @[WritebackQueue.scala 49:28]
  wire  serializer_io_out_ready; // @[WritebackQueue.scala 49:28]
  wire  serializer_io_out_valid; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_out_bits_0; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_out_bits_1; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_out_bits_2; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_out_bits_3; // @[WritebackQueue.scala 49:28]
  wire  serializer_io_fireAll; // @[WritebackQueue.scala 49:28]
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] reqReg_addr; // @[Reg.scala 19:16]
  reg [18:0] reqReg_dirtyTag; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_0; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_1; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_2; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_3; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire [18:0] _GEN_1 = _reqReg_T ? io_req_bits_dirtyTag : reqReg_dirtyTag; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_2 = _reqReg_T ? io_req_bits_data_0 : reqReg_data_0; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_3 = _reqReg_T ? io_req_bits_data_1 : reqReg_data_1; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_4 = _reqReg_T ? io_req_bits_data_2 : reqReg_data_2; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_5 = _reqReg_T ? io_req_bits_data_3 : reqReg_data_3; // @[Reg.scala 19:16 20:{18,22}]
  wire [18:0] req_dirtyTag = _reqReg_T ? io_req_bits_dirtyTag : reqReg_dirtyTag; // @[WritebackQueue.scala 43:18]
  reg  reqValidReg; // @[Reg.scala 19:16]
  wire  _GEN_6 = _reqReg_T | reqValidReg; // @[Reg.scala 19:16 20:{18,22}]
  wire [127:0] _T = {_GEN_5,_GEN_4,_GEN_3,_GEN_2}; // @[WritebackQueue.scala 51:47]
  reg [1:0] state; // @[WritebackQueue.scala 53:24]
  wire  _io_req_ready_T = state == 2'h0; // @[WritebackQueue.scala 56:27]
  wire  _GEN_8 = _io_req_ready_T & _reqReg_T; // @[WritebackQueue.scala 58:27 54:29]
  wire [1:0] _GEN_9 = serializer_io_fireAll ? 2'h2 : 2'h1; // @[WritebackQueue.scala 66:19 67:37 68:23]
  wire  _GEN_10 = serializer_io_fireAll ? 1'h0 : _GEN_6; // @[WritebackQueue.scala 67:37 70:25]
  wire  _GEN_12 = state == 2'h1 ? _GEN_10 : _GEN_6; // @[WritebackQueue.scala 65:34]
  wire  _T_8 = state == 2'h2; // @[WritebackQueue.scala 74:16]
  wire  _T_9 = io_tlbus_resp_ready & io_tlbus_resp_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_13 = io_resp_valid ? 2'h0 : 2'h3; // @[WritebackQueue.scala 77:23 79:32 80:27]
  wire  _T_11 = state == 2'h3; // @[WritebackQueue.scala 85:16]
  wire [63:0] io_tlbus_req_bits_data_lo = {serializer_io_out_bits_1,serializer_io_out_bits_0}; // @[WritebackQueue.scala 103:54]
  wire [63:0] io_tlbus_req_bits_data_hi = {serializer_io_out_bits_3,serializer_io_out_bits_2}; // @[WritebackQueue.scala 103:54]
  wire [8:0] dirtySet = _GEN_0[12:4]; // @[Parameters.scala 50:11]
  wire [31:0] writebackAddr = {_GEN_1,dirtySet,4'h0}; // @[Cat.scala 33:92]
  wire [32:0] _io_tlbus_req_bits_address_T_1 = {{1'd0}, writebackAddr}; // @[WritebackQueue.scala 110:49]
  TLSerializer serializer ( // @[WritebackQueue.scala 49:28]
    .io_in_valid(serializer_io_in_valid),
    .io_in_bits_0_0(serializer_io_in_bits_0_0),
    .io_in_bits_0_1(serializer_io_in_bits_0_1),
    .io_in_bits_0_2(serializer_io_in_bits_0_2),
    .io_in_bits_0_3(serializer_io_in_bits_0_3),
    .io_out_ready(serializer_io_out_ready),
    .io_out_valid(serializer_io_out_valid),
    .io_out_bits_0(serializer_io_out_bits_0),
    .io_out_bits_1(serializer_io_out_bits_1),
    .io_out_bits_2(serializer_io_out_bits_2),
    .io_out_bits_3(serializer_io_out_bits_3),
    .io_fireAll(serializer_io_fireAll)
  );
  assign io_req_ready = state == 2'h0; // @[WritebackQueue.scala 56:27]
  assign io_resp_valid = _T_11 | _T_9 & _T_8; // @[WritebackQueue.scala 96:38]
  assign io_tlbus_req_valid = serializer_io_out_valid; // @[WritebackQueue.scala 101:24]
  assign io_tlbus_req_bits_address = _io_tlbus_req_bits_address_T_1[31:0]; // @[WritebackQueue.scala 110:49]
  assign io_tlbus_req_bits_data = {io_tlbus_req_bits_data_hi,io_tlbus_req_bits_data_lo}; // @[WritebackQueue.scala 103:54]
  assign io_tlbus_resp_ready = 1'h1; // @[WritebackQueue.scala 98:25]
  assign serializer_io_in_valid = _reqReg_T | reqValidReg; // @[WritebackQueue.scala 45:23]
  assign serializer_io_in_bits_0_0 = _T[31:0]; // @[WritebackQueue.scala 51:47]
  assign serializer_io_in_bits_0_1 = _T[63:32]; // @[WritebackQueue.scala 51:47]
  assign serializer_io_in_bits_0_2 = _T[95:64]; // @[WritebackQueue.scala 51:47]
  assign serializer_io_in_bits_0_3 = _T[127:96]; // @[WritebackQueue.scala 51:47]
  assign serializer_io_out_ready = io_tlbus_req_ready; // @[WritebackQueue.scala 100:29]
  always @(posedge clock) begin
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_addr <= io_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_dirtyTag <= io_req_bits_dirtyTag; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_0 <= io_req_bits_data_0; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_1 <= io_req_bits_data_1; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_2 <= io_req_bits_data_2; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_3 <= io_req_bits_data_3; // @[Reg.scala 20:22]
    end
    if (state == 2'h3) begin // @[WritebackQueue.scala 85:27]
      if (io_resp_valid) begin // @[WritebackQueue.scala 87:28]
        reqValidReg <= 1'h0; // @[WritebackQueue.scala 90:25]
      end else begin
        reqValidReg <= _GEN_12;
      end
    end else begin
      reqValidReg <= _GEN_12;
    end
    if (reset) begin // @[WritebackQueue.scala 53:24]
      state <= 2'h0; // @[WritebackQueue.scala 53:24]
    end else if (state == 2'h3) begin // @[WritebackQueue.scala 85:27]
      state <= _GEN_13;
    end else if (state == 2'h2) begin // @[WritebackQueue.scala 74:32]
      if (_T_9) begin // @[WritebackQueue.scala 76:34]
        state <= _GEN_13;
      end else begin
        state <= 2'h2; // @[WritebackQueue.scala 75:19]
      end
    end else if (state == 2'h1) begin // @[WritebackQueue.scala 65:34]
      state <= _GEN_9;
    end else begin
      state <= {{1'd0}, _GEN_8};
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reqReg_addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reqReg_dirtyTag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  reqReg_data_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reqReg_data_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reqReg_data_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reqReg_data_3 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reqValidReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BankRAM_2P_80(
  input         clock,
  input         reset,
  input  [8:0]  io_r_addr,
  output [31:0] io_r_data,
  input         io_w_en,
  input  [8:0]  io_w_addr,
  input  [31:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:511]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_129_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_130_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_131_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_132_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_133_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_134_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_135_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_136_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_137_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_138_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_139_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_140_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_141_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_142_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_143_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_144_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_145_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_146_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_147_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_148_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_149_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_150_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_151_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_152_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_153_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_154_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_155_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_156_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_157_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_158_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_159_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_160_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_161_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_162_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_163_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_164_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_165_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_166_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_167_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_168_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_169_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_170_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_171_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_172_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_173_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_174_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_175_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_176_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_177_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_178_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_179_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_180_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_181_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_182_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_183_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_184_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_185_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_186_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_187_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_188_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_189_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_190_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_191_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_192_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_193_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_194_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_195_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_196_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_197_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_198_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_199_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_200_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_201_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_202_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_203_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_204_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_205_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_206_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_207_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_208_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_209_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_210_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_211_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_212_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_213_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_214_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_215_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_216_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_217_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_218_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_219_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_220_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_221_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_222_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_223_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_224_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_225_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_226_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_227_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_228_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_229_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_230_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_231_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_232_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_233_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_234_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_235_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_236_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_237_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_238_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_239_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_240_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_241_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_242_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_243_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_244_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_245_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_246_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_247_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_248_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_249_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_250_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_251_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_252_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_253_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_254_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_255_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_256_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_257_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_257_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_257_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_257_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_258_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_258_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_258_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_258_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_259_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_259_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_259_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_259_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_260_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_260_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_260_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_260_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_261_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_261_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_261_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_261_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_262_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_262_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_262_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_262_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_263_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_263_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_263_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_263_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_264_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_264_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_264_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_264_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_265_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_265_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_265_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_265_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_266_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_266_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_266_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_266_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_267_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_267_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_267_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_267_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_268_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_268_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_268_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_268_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_269_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_269_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_269_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_269_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_270_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_270_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_270_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_270_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_271_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_271_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_271_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_271_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_272_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_272_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_272_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_272_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_273_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_273_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_273_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_273_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_274_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_274_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_274_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_274_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_275_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_275_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_275_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_275_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_276_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_276_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_276_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_276_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_277_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_277_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_277_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_277_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_278_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_278_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_278_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_278_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_279_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_279_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_279_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_279_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_280_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_280_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_280_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_280_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_281_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_281_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_281_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_281_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_282_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_282_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_282_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_282_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_283_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_283_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_283_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_283_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_284_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_284_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_284_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_284_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_285_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_285_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_285_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_285_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_286_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_286_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_286_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_286_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_287_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_287_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_287_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_287_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_288_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_288_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_288_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_288_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_289_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_289_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_289_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_289_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_290_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_290_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_290_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_290_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_291_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_291_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_291_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_291_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_292_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_292_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_292_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_292_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_293_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_293_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_293_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_293_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_294_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_294_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_294_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_294_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_295_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_295_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_295_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_295_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_296_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_296_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_296_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_296_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_297_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_297_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_297_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_297_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_298_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_298_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_298_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_298_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_299_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_299_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_299_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_299_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_300_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_300_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_300_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_300_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_301_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_301_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_301_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_301_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_302_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_302_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_302_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_302_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_303_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_303_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_303_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_303_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_304_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_304_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_304_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_304_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_305_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_305_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_305_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_305_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_306_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_306_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_306_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_306_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_307_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_307_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_307_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_307_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_308_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_308_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_308_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_308_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_309_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_309_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_309_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_309_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_310_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_310_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_310_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_310_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_311_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_311_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_311_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_311_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_312_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_312_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_312_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_312_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_313_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_313_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_313_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_313_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_314_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_314_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_314_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_314_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_315_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_315_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_315_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_315_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_316_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_316_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_316_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_316_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_317_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_317_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_317_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_317_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_318_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_318_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_318_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_318_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_319_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_319_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_319_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_319_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_320_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_320_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_320_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_320_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_321_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_321_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_321_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_321_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_322_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_322_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_322_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_322_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_323_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_323_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_323_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_323_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_324_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_324_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_324_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_324_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_325_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_325_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_325_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_325_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_326_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_326_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_326_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_326_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_327_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_327_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_327_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_327_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_328_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_328_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_328_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_328_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_329_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_329_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_329_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_329_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_330_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_330_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_330_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_330_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_331_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_331_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_331_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_331_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_332_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_332_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_332_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_332_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_333_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_333_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_333_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_333_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_334_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_334_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_334_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_334_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_335_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_335_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_335_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_335_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_336_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_336_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_336_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_336_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_337_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_337_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_337_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_337_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_338_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_338_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_338_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_338_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_339_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_339_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_339_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_339_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_340_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_340_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_340_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_340_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_341_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_341_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_341_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_341_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_342_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_342_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_342_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_342_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_343_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_343_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_343_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_343_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_344_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_344_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_344_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_344_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_345_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_345_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_345_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_345_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_346_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_346_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_346_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_346_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_347_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_347_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_347_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_347_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_348_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_348_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_348_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_348_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_349_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_349_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_349_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_349_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_350_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_350_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_350_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_350_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_351_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_351_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_351_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_351_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_352_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_352_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_352_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_352_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_353_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_353_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_353_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_353_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_354_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_354_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_354_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_354_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_355_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_355_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_355_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_355_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_356_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_356_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_356_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_356_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_357_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_357_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_357_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_357_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_358_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_358_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_358_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_358_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_359_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_359_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_359_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_359_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_360_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_360_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_360_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_360_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_361_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_361_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_361_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_361_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_362_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_362_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_362_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_362_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_363_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_363_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_363_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_363_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_364_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_364_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_364_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_364_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_365_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_365_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_365_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_365_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_366_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_366_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_366_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_366_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_367_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_367_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_367_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_367_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_368_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_368_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_368_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_368_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_369_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_369_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_369_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_369_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_370_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_370_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_370_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_370_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_371_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_371_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_371_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_371_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_372_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_372_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_372_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_372_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_373_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_373_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_373_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_373_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_374_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_374_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_374_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_374_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_375_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_375_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_375_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_375_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_376_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_376_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_376_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_376_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_377_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_377_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_377_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_377_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_378_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_378_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_378_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_378_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_379_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_379_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_379_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_379_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_380_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_380_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_380_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_380_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_381_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_381_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_381_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_381_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_382_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_382_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_382_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_382_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_383_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_383_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_383_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_383_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_384_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_384_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_384_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_384_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_385_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_385_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_385_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_385_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_386_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_386_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_386_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_386_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_387_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_387_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_387_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_387_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_388_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_388_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_388_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_388_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_389_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_389_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_389_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_389_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_390_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_390_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_390_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_390_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_391_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_391_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_391_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_391_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_392_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_392_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_392_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_392_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_393_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_393_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_393_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_393_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_394_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_394_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_394_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_394_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_395_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_395_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_395_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_395_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_396_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_396_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_396_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_396_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_397_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_397_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_397_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_397_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_398_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_398_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_398_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_398_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_399_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_399_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_399_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_399_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_400_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_400_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_400_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_400_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_401_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_401_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_401_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_401_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_402_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_402_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_402_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_402_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_403_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_403_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_403_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_403_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_404_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_404_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_404_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_404_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_405_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_405_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_405_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_405_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_406_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_406_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_406_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_406_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_407_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_407_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_407_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_407_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_408_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_408_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_408_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_408_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_409_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_409_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_409_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_409_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_410_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_410_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_410_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_410_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_411_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_411_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_411_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_411_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_412_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_412_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_412_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_412_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_413_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_413_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_413_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_413_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_414_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_414_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_414_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_414_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_415_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_415_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_415_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_415_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_416_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_416_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_416_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_416_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_417_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_417_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_417_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_417_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_418_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_418_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_418_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_418_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_419_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_419_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_419_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_419_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_420_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_420_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_420_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_420_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_421_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_421_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_421_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_421_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_422_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_422_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_422_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_422_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_423_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_423_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_423_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_423_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_424_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_424_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_424_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_424_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_425_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_425_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_425_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_425_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_426_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_426_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_426_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_426_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_427_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_427_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_427_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_427_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_428_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_428_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_428_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_428_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_429_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_429_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_429_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_429_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_430_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_430_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_430_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_430_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_431_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_431_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_431_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_431_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_432_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_432_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_432_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_432_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_433_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_433_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_433_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_433_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_434_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_434_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_434_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_434_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_435_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_435_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_435_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_435_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_436_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_436_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_436_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_436_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_437_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_437_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_437_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_437_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_438_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_438_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_438_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_438_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_439_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_439_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_439_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_439_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_440_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_440_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_440_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_440_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_441_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_441_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_441_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_441_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_442_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_442_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_442_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_442_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_443_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_443_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_443_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_443_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_444_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_444_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_444_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_444_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_445_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_445_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_445_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_445_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_446_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_446_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_446_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_446_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_447_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_447_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_447_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_447_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_448_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_448_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_448_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_448_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_449_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_449_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_449_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_449_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_450_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_450_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_450_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_450_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_451_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_451_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_451_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_451_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_452_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_452_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_452_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_452_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_453_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_453_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_453_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_453_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_454_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_454_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_454_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_454_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_455_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_455_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_455_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_455_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_456_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_456_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_456_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_456_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_457_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_457_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_457_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_457_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_458_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_458_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_458_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_458_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_459_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_459_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_459_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_459_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_460_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_460_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_460_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_460_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_461_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_461_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_461_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_461_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_462_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_462_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_462_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_462_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_463_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_463_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_463_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_463_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_464_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_464_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_464_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_464_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_465_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_465_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_465_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_465_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_466_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_466_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_466_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_466_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_467_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_467_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_467_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_467_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_468_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_468_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_468_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_468_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_469_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_469_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_469_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_469_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_470_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_470_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_470_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_470_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_471_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_471_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_471_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_471_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_472_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_472_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_472_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_472_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_473_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_473_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_473_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_473_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_474_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_474_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_474_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_474_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_475_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_475_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_475_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_475_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_476_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_476_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_476_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_476_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_477_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_477_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_477_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_477_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_478_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_478_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_478_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_478_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_479_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_479_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_479_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_479_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_480_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_480_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_480_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_480_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_481_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_481_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_481_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_481_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_482_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_482_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_482_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_482_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_483_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_483_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_483_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_483_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_484_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_484_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_484_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_484_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_485_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_485_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_485_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_485_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_486_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_486_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_486_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_486_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_487_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_487_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_487_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_487_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_488_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_488_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_488_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_488_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_489_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_489_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_489_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_489_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_490_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_490_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_490_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_490_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_491_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_491_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_491_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_491_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_492_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_492_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_492_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_492_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_493_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_493_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_493_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_493_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_494_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_494_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_494_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_494_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_495_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_495_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_495_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_495_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_496_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_496_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_496_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_496_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_497_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_497_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_497_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_497_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_498_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_498_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_498_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_498_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_499_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_499_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_499_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_499_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_500_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_500_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_500_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_500_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_501_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_501_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_501_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_501_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_502_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_502_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_502_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_502_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_503_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_503_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_503_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_503_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_504_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_504_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_504_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_504_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_505_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_505_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_505_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_505_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_506_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_506_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_506_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_506_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_507_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_507_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_507_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_507_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_508_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_508_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_508_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_508_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_509_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_509_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_509_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_509_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_510_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_510_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_510_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_510_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_511_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_511_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_511_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_511_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_512_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_512_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_512_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_512_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [8:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 32'h0;
  assign mem_MPORT_addr = 9'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 32'h0;
  assign mem_MPORT_1_addr = 9'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 32'h0;
  assign mem_MPORT_2_addr = 9'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 32'h0;
  assign mem_MPORT_3_addr = 9'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 32'h0;
  assign mem_MPORT_4_addr = 9'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 32'h0;
  assign mem_MPORT_5_addr = 9'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 32'h0;
  assign mem_MPORT_6_addr = 9'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 32'h0;
  assign mem_MPORT_7_addr = 9'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 32'h0;
  assign mem_MPORT_8_addr = 9'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 32'h0;
  assign mem_MPORT_9_addr = 9'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 32'h0;
  assign mem_MPORT_10_addr = 9'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 32'h0;
  assign mem_MPORT_11_addr = 9'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 32'h0;
  assign mem_MPORT_12_addr = 9'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 32'h0;
  assign mem_MPORT_13_addr = 9'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 32'h0;
  assign mem_MPORT_14_addr = 9'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 32'h0;
  assign mem_MPORT_15_addr = 9'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 32'h0;
  assign mem_MPORT_16_addr = 9'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 32'h0;
  assign mem_MPORT_17_addr = 9'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 32'h0;
  assign mem_MPORT_18_addr = 9'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 32'h0;
  assign mem_MPORT_19_addr = 9'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 32'h0;
  assign mem_MPORT_20_addr = 9'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 32'h0;
  assign mem_MPORT_21_addr = 9'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 32'h0;
  assign mem_MPORT_22_addr = 9'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 32'h0;
  assign mem_MPORT_23_addr = 9'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 32'h0;
  assign mem_MPORT_24_addr = 9'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 32'h0;
  assign mem_MPORT_25_addr = 9'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 32'h0;
  assign mem_MPORT_26_addr = 9'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 32'h0;
  assign mem_MPORT_27_addr = 9'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 32'h0;
  assign mem_MPORT_28_addr = 9'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 32'h0;
  assign mem_MPORT_29_addr = 9'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 32'h0;
  assign mem_MPORT_30_addr = 9'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 32'h0;
  assign mem_MPORT_31_addr = 9'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 32'h0;
  assign mem_MPORT_32_addr = 9'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 32'h0;
  assign mem_MPORT_33_addr = 9'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 32'h0;
  assign mem_MPORT_34_addr = 9'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 32'h0;
  assign mem_MPORT_35_addr = 9'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 32'h0;
  assign mem_MPORT_36_addr = 9'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 32'h0;
  assign mem_MPORT_37_addr = 9'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 32'h0;
  assign mem_MPORT_38_addr = 9'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 32'h0;
  assign mem_MPORT_39_addr = 9'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 32'h0;
  assign mem_MPORT_40_addr = 9'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 32'h0;
  assign mem_MPORT_41_addr = 9'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 32'h0;
  assign mem_MPORT_42_addr = 9'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 32'h0;
  assign mem_MPORT_43_addr = 9'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 32'h0;
  assign mem_MPORT_44_addr = 9'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 32'h0;
  assign mem_MPORT_45_addr = 9'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 32'h0;
  assign mem_MPORT_46_addr = 9'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 32'h0;
  assign mem_MPORT_47_addr = 9'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 32'h0;
  assign mem_MPORT_48_addr = 9'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 32'h0;
  assign mem_MPORT_49_addr = 9'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 32'h0;
  assign mem_MPORT_50_addr = 9'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 32'h0;
  assign mem_MPORT_51_addr = 9'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 32'h0;
  assign mem_MPORT_52_addr = 9'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 32'h0;
  assign mem_MPORT_53_addr = 9'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 32'h0;
  assign mem_MPORT_54_addr = 9'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 32'h0;
  assign mem_MPORT_55_addr = 9'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 32'h0;
  assign mem_MPORT_56_addr = 9'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 32'h0;
  assign mem_MPORT_57_addr = 9'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 32'h0;
  assign mem_MPORT_58_addr = 9'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 32'h0;
  assign mem_MPORT_59_addr = 9'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 32'h0;
  assign mem_MPORT_60_addr = 9'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 32'h0;
  assign mem_MPORT_61_addr = 9'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 32'h0;
  assign mem_MPORT_62_addr = 9'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 32'h0;
  assign mem_MPORT_63_addr = 9'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 32'h0;
  assign mem_MPORT_64_addr = 9'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 32'h0;
  assign mem_MPORT_65_addr = 9'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 32'h0;
  assign mem_MPORT_66_addr = 9'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 32'h0;
  assign mem_MPORT_67_addr = 9'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 32'h0;
  assign mem_MPORT_68_addr = 9'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 32'h0;
  assign mem_MPORT_69_addr = 9'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 32'h0;
  assign mem_MPORT_70_addr = 9'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 32'h0;
  assign mem_MPORT_71_addr = 9'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 32'h0;
  assign mem_MPORT_72_addr = 9'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 32'h0;
  assign mem_MPORT_73_addr = 9'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 32'h0;
  assign mem_MPORT_74_addr = 9'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 32'h0;
  assign mem_MPORT_75_addr = 9'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 32'h0;
  assign mem_MPORT_76_addr = 9'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 32'h0;
  assign mem_MPORT_77_addr = 9'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 32'h0;
  assign mem_MPORT_78_addr = 9'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 32'h0;
  assign mem_MPORT_79_addr = 9'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 32'h0;
  assign mem_MPORT_80_addr = 9'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 32'h0;
  assign mem_MPORT_81_addr = 9'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 32'h0;
  assign mem_MPORT_82_addr = 9'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 32'h0;
  assign mem_MPORT_83_addr = 9'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 32'h0;
  assign mem_MPORT_84_addr = 9'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 32'h0;
  assign mem_MPORT_85_addr = 9'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 32'h0;
  assign mem_MPORT_86_addr = 9'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 32'h0;
  assign mem_MPORT_87_addr = 9'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 32'h0;
  assign mem_MPORT_88_addr = 9'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 32'h0;
  assign mem_MPORT_89_addr = 9'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 32'h0;
  assign mem_MPORT_90_addr = 9'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 32'h0;
  assign mem_MPORT_91_addr = 9'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 32'h0;
  assign mem_MPORT_92_addr = 9'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 32'h0;
  assign mem_MPORT_93_addr = 9'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 32'h0;
  assign mem_MPORT_94_addr = 9'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 32'h0;
  assign mem_MPORT_95_addr = 9'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 32'h0;
  assign mem_MPORT_96_addr = 9'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 32'h0;
  assign mem_MPORT_97_addr = 9'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 32'h0;
  assign mem_MPORT_98_addr = 9'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 32'h0;
  assign mem_MPORT_99_addr = 9'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 32'h0;
  assign mem_MPORT_100_addr = 9'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 32'h0;
  assign mem_MPORT_101_addr = 9'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 32'h0;
  assign mem_MPORT_102_addr = 9'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 32'h0;
  assign mem_MPORT_103_addr = 9'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 32'h0;
  assign mem_MPORT_104_addr = 9'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 32'h0;
  assign mem_MPORT_105_addr = 9'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 32'h0;
  assign mem_MPORT_106_addr = 9'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 32'h0;
  assign mem_MPORT_107_addr = 9'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 32'h0;
  assign mem_MPORT_108_addr = 9'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 32'h0;
  assign mem_MPORT_109_addr = 9'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 32'h0;
  assign mem_MPORT_110_addr = 9'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 32'h0;
  assign mem_MPORT_111_addr = 9'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 32'h0;
  assign mem_MPORT_112_addr = 9'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 32'h0;
  assign mem_MPORT_113_addr = 9'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 32'h0;
  assign mem_MPORT_114_addr = 9'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 32'h0;
  assign mem_MPORT_115_addr = 9'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 32'h0;
  assign mem_MPORT_116_addr = 9'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 32'h0;
  assign mem_MPORT_117_addr = 9'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 32'h0;
  assign mem_MPORT_118_addr = 9'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 32'h0;
  assign mem_MPORT_119_addr = 9'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 32'h0;
  assign mem_MPORT_120_addr = 9'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 32'h0;
  assign mem_MPORT_121_addr = 9'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 32'h0;
  assign mem_MPORT_122_addr = 9'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 32'h0;
  assign mem_MPORT_123_addr = 9'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 32'h0;
  assign mem_MPORT_124_addr = 9'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 32'h0;
  assign mem_MPORT_125_addr = 9'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 32'h0;
  assign mem_MPORT_126_addr = 9'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 32'h0;
  assign mem_MPORT_127_addr = 9'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 32'h0;
  assign mem_MPORT_128_addr = 9'h80;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = reset;
  assign mem_MPORT_129_data = 32'h0;
  assign mem_MPORT_129_addr = 9'h81;
  assign mem_MPORT_129_mask = 1'h1;
  assign mem_MPORT_129_en = reset;
  assign mem_MPORT_130_data = 32'h0;
  assign mem_MPORT_130_addr = 9'h82;
  assign mem_MPORT_130_mask = 1'h1;
  assign mem_MPORT_130_en = reset;
  assign mem_MPORT_131_data = 32'h0;
  assign mem_MPORT_131_addr = 9'h83;
  assign mem_MPORT_131_mask = 1'h1;
  assign mem_MPORT_131_en = reset;
  assign mem_MPORT_132_data = 32'h0;
  assign mem_MPORT_132_addr = 9'h84;
  assign mem_MPORT_132_mask = 1'h1;
  assign mem_MPORT_132_en = reset;
  assign mem_MPORT_133_data = 32'h0;
  assign mem_MPORT_133_addr = 9'h85;
  assign mem_MPORT_133_mask = 1'h1;
  assign mem_MPORT_133_en = reset;
  assign mem_MPORT_134_data = 32'h0;
  assign mem_MPORT_134_addr = 9'h86;
  assign mem_MPORT_134_mask = 1'h1;
  assign mem_MPORT_134_en = reset;
  assign mem_MPORT_135_data = 32'h0;
  assign mem_MPORT_135_addr = 9'h87;
  assign mem_MPORT_135_mask = 1'h1;
  assign mem_MPORT_135_en = reset;
  assign mem_MPORT_136_data = 32'h0;
  assign mem_MPORT_136_addr = 9'h88;
  assign mem_MPORT_136_mask = 1'h1;
  assign mem_MPORT_136_en = reset;
  assign mem_MPORT_137_data = 32'h0;
  assign mem_MPORT_137_addr = 9'h89;
  assign mem_MPORT_137_mask = 1'h1;
  assign mem_MPORT_137_en = reset;
  assign mem_MPORT_138_data = 32'h0;
  assign mem_MPORT_138_addr = 9'h8a;
  assign mem_MPORT_138_mask = 1'h1;
  assign mem_MPORT_138_en = reset;
  assign mem_MPORT_139_data = 32'h0;
  assign mem_MPORT_139_addr = 9'h8b;
  assign mem_MPORT_139_mask = 1'h1;
  assign mem_MPORT_139_en = reset;
  assign mem_MPORT_140_data = 32'h0;
  assign mem_MPORT_140_addr = 9'h8c;
  assign mem_MPORT_140_mask = 1'h1;
  assign mem_MPORT_140_en = reset;
  assign mem_MPORT_141_data = 32'h0;
  assign mem_MPORT_141_addr = 9'h8d;
  assign mem_MPORT_141_mask = 1'h1;
  assign mem_MPORT_141_en = reset;
  assign mem_MPORT_142_data = 32'h0;
  assign mem_MPORT_142_addr = 9'h8e;
  assign mem_MPORT_142_mask = 1'h1;
  assign mem_MPORT_142_en = reset;
  assign mem_MPORT_143_data = 32'h0;
  assign mem_MPORT_143_addr = 9'h8f;
  assign mem_MPORT_143_mask = 1'h1;
  assign mem_MPORT_143_en = reset;
  assign mem_MPORT_144_data = 32'h0;
  assign mem_MPORT_144_addr = 9'h90;
  assign mem_MPORT_144_mask = 1'h1;
  assign mem_MPORT_144_en = reset;
  assign mem_MPORT_145_data = 32'h0;
  assign mem_MPORT_145_addr = 9'h91;
  assign mem_MPORT_145_mask = 1'h1;
  assign mem_MPORT_145_en = reset;
  assign mem_MPORT_146_data = 32'h0;
  assign mem_MPORT_146_addr = 9'h92;
  assign mem_MPORT_146_mask = 1'h1;
  assign mem_MPORT_146_en = reset;
  assign mem_MPORT_147_data = 32'h0;
  assign mem_MPORT_147_addr = 9'h93;
  assign mem_MPORT_147_mask = 1'h1;
  assign mem_MPORT_147_en = reset;
  assign mem_MPORT_148_data = 32'h0;
  assign mem_MPORT_148_addr = 9'h94;
  assign mem_MPORT_148_mask = 1'h1;
  assign mem_MPORT_148_en = reset;
  assign mem_MPORT_149_data = 32'h0;
  assign mem_MPORT_149_addr = 9'h95;
  assign mem_MPORT_149_mask = 1'h1;
  assign mem_MPORT_149_en = reset;
  assign mem_MPORT_150_data = 32'h0;
  assign mem_MPORT_150_addr = 9'h96;
  assign mem_MPORT_150_mask = 1'h1;
  assign mem_MPORT_150_en = reset;
  assign mem_MPORT_151_data = 32'h0;
  assign mem_MPORT_151_addr = 9'h97;
  assign mem_MPORT_151_mask = 1'h1;
  assign mem_MPORT_151_en = reset;
  assign mem_MPORT_152_data = 32'h0;
  assign mem_MPORT_152_addr = 9'h98;
  assign mem_MPORT_152_mask = 1'h1;
  assign mem_MPORT_152_en = reset;
  assign mem_MPORT_153_data = 32'h0;
  assign mem_MPORT_153_addr = 9'h99;
  assign mem_MPORT_153_mask = 1'h1;
  assign mem_MPORT_153_en = reset;
  assign mem_MPORT_154_data = 32'h0;
  assign mem_MPORT_154_addr = 9'h9a;
  assign mem_MPORT_154_mask = 1'h1;
  assign mem_MPORT_154_en = reset;
  assign mem_MPORT_155_data = 32'h0;
  assign mem_MPORT_155_addr = 9'h9b;
  assign mem_MPORT_155_mask = 1'h1;
  assign mem_MPORT_155_en = reset;
  assign mem_MPORT_156_data = 32'h0;
  assign mem_MPORT_156_addr = 9'h9c;
  assign mem_MPORT_156_mask = 1'h1;
  assign mem_MPORT_156_en = reset;
  assign mem_MPORT_157_data = 32'h0;
  assign mem_MPORT_157_addr = 9'h9d;
  assign mem_MPORT_157_mask = 1'h1;
  assign mem_MPORT_157_en = reset;
  assign mem_MPORT_158_data = 32'h0;
  assign mem_MPORT_158_addr = 9'h9e;
  assign mem_MPORT_158_mask = 1'h1;
  assign mem_MPORT_158_en = reset;
  assign mem_MPORT_159_data = 32'h0;
  assign mem_MPORT_159_addr = 9'h9f;
  assign mem_MPORT_159_mask = 1'h1;
  assign mem_MPORT_159_en = reset;
  assign mem_MPORT_160_data = 32'h0;
  assign mem_MPORT_160_addr = 9'ha0;
  assign mem_MPORT_160_mask = 1'h1;
  assign mem_MPORT_160_en = reset;
  assign mem_MPORT_161_data = 32'h0;
  assign mem_MPORT_161_addr = 9'ha1;
  assign mem_MPORT_161_mask = 1'h1;
  assign mem_MPORT_161_en = reset;
  assign mem_MPORT_162_data = 32'h0;
  assign mem_MPORT_162_addr = 9'ha2;
  assign mem_MPORT_162_mask = 1'h1;
  assign mem_MPORT_162_en = reset;
  assign mem_MPORT_163_data = 32'h0;
  assign mem_MPORT_163_addr = 9'ha3;
  assign mem_MPORT_163_mask = 1'h1;
  assign mem_MPORT_163_en = reset;
  assign mem_MPORT_164_data = 32'h0;
  assign mem_MPORT_164_addr = 9'ha4;
  assign mem_MPORT_164_mask = 1'h1;
  assign mem_MPORT_164_en = reset;
  assign mem_MPORT_165_data = 32'h0;
  assign mem_MPORT_165_addr = 9'ha5;
  assign mem_MPORT_165_mask = 1'h1;
  assign mem_MPORT_165_en = reset;
  assign mem_MPORT_166_data = 32'h0;
  assign mem_MPORT_166_addr = 9'ha6;
  assign mem_MPORT_166_mask = 1'h1;
  assign mem_MPORT_166_en = reset;
  assign mem_MPORT_167_data = 32'h0;
  assign mem_MPORT_167_addr = 9'ha7;
  assign mem_MPORT_167_mask = 1'h1;
  assign mem_MPORT_167_en = reset;
  assign mem_MPORT_168_data = 32'h0;
  assign mem_MPORT_168_addr = 9'ha8;
  assign mem_MPORT_168_mask = 1'h1;
  assign mem_MPORT_168_en = reset;
  assign mem_MPORT_169_data = 32'h0;
  assign mem_MPORT_169_addr = 9'ha9;
  assign mem_MPORT_169_mask = 1'h1;
  assign mem_MPORT_169_en = reset;
  assign mem_MPORT_170_data = 32'h0;
  assign mem_MPORT_170_addr = 9'haa;
  assign mem_MPORT_170_mask = 1'h1;
  assign mem_MPORT_170_en = reset;
  assign mem_MPORT_171_data = 32'h0;
  assign mem_MPORT_171_addr = 9'hab;
  assign mem_MPORT_171_mask = 1'h1;
  assign mem_MPORT_171_en = reset;
  assign mem_MPORT_172_data = 32'h0;
  assign mem_MPORT_172_addr = 9'hac;
  assign mem_MPORT_172_mask = 1'h1;
  assign mem_MPORT_172_en = reset;
  assign mem_MPORT_173_data = 32'h0;
  assign mem_MPORT_173_addr = 9'had;
  assign mem_MPORT_173_mask = 1'h1;
  assign mem_MPORT_173_en = reset;
  assign mem_MPORT_174_data = 32'h0;
  assign mem_MPORT_174_addr = 9'hae;
  assign mem_MPORT_174_mask = 1'h1;
  assign mem_MPORT_174_en = reset;
  assign mem_MPORT_175_data = 32'h0;
  assign mem_MPORT_175_addr = 9'haf;
  assign mem_MPORT_175_mask = 1'h1;
  assign mem_MPORT_175_en = reset;
  assign mem_MPORT_176_data = 32'h0;
  assign mem_MPORT_176_addr = 9'hb0;
  assign mem_MPORT_176_mask = 1'h1;
  assign mem_MPORT_176_en = reset;
  assign mem_MPORT_177_data = 32'h0;
  assign mem_MPORT_177_addr = 9'hb1;
  assign mem_MPORT_177_mask = 1'h1;
  assign mem_MPORT_177_en = reset;
  assign mem_MPORT_178_data = 32'h0;
  assign mem_MPORT_178_addr = 9'hb2;
  assign mem_MPORT_178_mask = 1'h1;
  assign mem_MPORT_178_en = reset;
  assign mem_MPORT_179_data = 32'h0;
  assign mem_MPORT_179_addr = 9'hb3;
  assign mem_MPORT_179_mask = 1'h1;
  assign mem_MPORT_179_en = reset;
  assign mem_MPORT_180_data = 32'h0;
  assign mem_MPORT_180_addr = 9'hb4;
  assign mem_MPORT_180_mask = 1'h1;
  assign mem_MPORT_180_en = reset;
  assign mem_MPORT_181_data = 32'h0;
  assign mem_MPORT_181_addr = 9'hb5;
  assign mem_MPORT_181_mask = 1'h1;
  assign mem_MPORT_181_en = reset;
  assign mem_MPORT_182_data = 32'h0;
  assign mem_MPORT_182_addr = 9'hb6;
  assign mem_MPORT_182_mask = 1'h1;
  assign mem_MPORT_182_en = reset;
  assign mem_MPORT_183_data = 32'h0;
  assign mem_MPORT_183_addr = 9'hb7;
  assign mem_MPORT_183_mask = 1'h1;
  assign mem_MPORT_183_en = reset;
  assign mem_MPORT_184_data = 32'h0;
  assign mem_MPORT_184_addr = 9'hb8;
  assign mem_MPORT_184_mask = 1'h1;
  assign mem_MPORT_184_en = reset;
  assign mem_MPORT_185_data = 32'h0;
  assign mem_MPORT_185_addr = 9'hb9;
  assign mem_MPORT_185_mask = 1'h1;
  assign mem_MPORT_185_en = reset;
  assign mem_MPORT_186_data = 32'h0;
  assign mem_MPORT_186_addr = 9'hba;
  assign mem_MPORT_186_mask = 1'h1;
  assign mem_MPORT_186_en = reset;
  assign mem_MPORT_187_data = 32'h0;
  assign mem_MPORT_187_addr = 9'hbb;
  assign mem_MPORT_187_mask = 1'h1;
  assign mem_MPORT_187_en = reset;
  assign mem_MPORT_188_data = 32'h0;
  assign mem_MPORT_188_addr = 9'hbc;
  assign mem_MPORT_188_mask = 1'h1;
  assign mem_MPORT_188_en = reset;
  assign mem_MPORT_189_data = 32'h0;
  assign mem_MPORT_189_addr = 9'hbd;
  assign mem_MPORT_189_mask = 1'h1;
  assign mem_MPORT_189_en = reset;
  assign mem_MPORT_190_data = 32'h0;
  assign mem_MPORT_190_addr = 9'hbe;
  assign mem_MPORT_190_mask = 1'h1;
  assign mem_MPORT_190_en = reset;
  assign mem_MPORT_191_data = 32'h0;
  assign mem_MPORT_191_addr = 9'hbf;
  assign mem_MPORT_191_mask = 1'h1;
  assign mem_MPORT_191_en = reset;
  assign mem_MPORT_192_data = 32'h0;
  assign mem_MPORT_192_addr = 9'hc0;
  assign mem_MPORT_192_mask = 1'h1;
  assign mem_MPORT_192_en = reset;
  assign mem_MPORT_193_data = 32'h0;
  assign mem_MPORT_193_addr = 9'hc1;
  assign mem_MPORT_193_mask = 1'h1;
  assign mem_MPORT_193_en = reset;
  assign mem_MPORT_194_data = 32'h0;
  assign mem_MPORT_194_addr = 9'hc2;
  assign mem_MPORT_194_mask = 1'h1;
  assign mem_MPORT_194_en = reset;
  assign mem_MPORT_195_data = 32'h0;
  assign mem_MPORT_195_addr = 9'hc3;
  assign mem_MPORT_195_mask = 1'h1;
  assign mem_MPORT_195_en = reset;
  assign mem_MPORT_196_data = 32'h0;
  assign mem_MPORT_196_addr = 9'hc4;
  assign mem_MPORT_196_mask = 1'h1;
  assign mem_MPORT_196_en = reset;
  assign mem_MPORT_197_data = 32'h0;
  assign mem_MPORT_197_addr = 9'hc5;
  assign mem_MPORT_197_mask = 1'h1;
  assign mem_MPORT_197_en = reset;
  assign mem_MPORT_198_data = 32'h0;
  assign mem_MPORT_198_addr = 9'hc6;
  assign mem_MPORT_198_mask = 1'h1;
  assign mem_MPORT_198_en = reset;
  assign mem_MPORT_199_data = 32'h0;
  assign mem_MPORT_199_addr = 9'hc7;
  assign mem_MPORT_199_mask = 1'h1;
  assign mem_MPORT_199_en = reset;
  assign mem_MPORT_200_data = 32'h0;
  assign mem_MPORT_200_addr = 9'hc8;
  assign mem_MPORT_200_mask = 1'h1;
  assign mem_MPORT_200_en = reset;
  assign mem_MPORT_201_data = 32'h0;
  assign mem_MPORT_201_addr = 9'hc9;
  assign mem_MPORT_201_mask = 1'h1;
  assign mem_MPORT_201_en = reset;
  assign mem_MPORT_202_data = 32'h0;
  assign mem_MPORT_202_addr = 9'hca;
  assign mem_MPORT_202_mask = 1'h1;
  assign mem_MPORT_202_en = reset;
  assign mem_MPORT_203_data = 32'h0;
  assign mem_MPORT_203_addr = 9'hcb;
  assign mem_MPORT_203_mask = 1'h1;
  assign mem_MPORT_203_en = reset;
  assign mem_MPORT_204_data = 32'h0;
  assign mem_MPORT_204_addr = 9'hcc;
  assign mem_MPORT_204_mask = 1'h1;
  assign mem_MPORT_204_en = reset;
  assign mem_MPORT_205_data = 32'h0;
  assign mem_MPORT_205_addr = 9'hcd;
  assign mem_MPORT_205_mask = 1'h1;
  assign mem_MPORT_205_en = reset;
  assign mem_MPORT_206_data = 32'h0;
  assign mem_MPORT_206_addr = 9'hce;
  assign mem_MPORT_206_mask = 1'h1;
  assign mem_MPORT_206_en = reset;
  assign mem_MPORT_207_data = 32'h0;
  assign mem_MPORT_207_addr = 9'hcf;
  assign mem_MPORT_207_mask = 1'h1;
  assign mem_MPORT_207_en = reset;
  assign mem_MPORT_208_data = 32'h0;
  assign mem_MPORT_208_addr = 9'hd0;
  assign mem_MPORT_208_mask = 1'h1;
  assign mem_MPORT_208_en = reset;
  assign mem_MPORT_209_data = 32'h0;
  assign mem_MPORT_209_addr = 9'hd1;
  assign mem_MPORT_209_mask = 1'h1;
  assign mem_MPORT_209_en = reset;
  assign mem_MPORT_210_data = 32'h0;
  assign mem_MPORT_210_addr = 9'hd2;
  assign mem_MPORT_210_mask = 1'h1;
  assign mem_MPORT_210_en = reset;
  assign mem_MPORT_211_data = 32'h0;
  assign mem_MPORT_211_addr = 9'hd3;
  assign mem_MPORT_211_mask = 1'h1;
  assign mem_MPORT_211_en = reset;
  assign mem_MPORT_212_data = 32'h0;
  assign mem_MPORT_212_addr = 9'hd4;
  assign mem_MPORT_212_mask = 1'h1;
  assign mem_MPORT_212_en = reset;
  assign mem_MPORT_213_data = 32'h0;
  assign mem_MPORT_213_addr = 9'hd5;
  assign mem_MPORT_213_mask = 1'h1;
  assign mem_MPORT_213_en = reset;
  assign mem_MPORT_214_data = 32'h0;
  assign mem_MPORT_214_addr = 9'hd6;
  assign mem_MPORT_214_mask = 1'h1;
  assign mem_MPORT_214_en = reset;
  assign mem_MPORT_215_data = 32'h0;
  assign mem_MPORT_215_addr = 9'hd7;
  assign mem_MPORT_215_mask = 1'h1;
  assign mem_MPORT_215_en = reset;
  assign mem_MPORT_216_data = 32'h0;
  assign mem_MPORT_216_addr = 9'hd8;
  assign mem_MPORT_216_mask = 1'h1;
  assign mem_MPORT_216_en = reset;
  assign mem_MPORT_217_data = 32'h0;
  assign mem_MPORT_217_addr = 9'hd9;
  assign mem_MPORT_217_mask = 1'h1;
  assign mem_MPORT_217_en = reset;
  assign mem_MPORT_218_data = 32'h0;
  assign mem_MPORT_218_addr = 9'hda;
  assign mem_MPORT_218_mask = 1'h1;
  assign mem_MPORT_218_en = reset;
  assign mem_MPORT_219_data = 32'h0;
  assign mem_MPORT_219_addr = 9'hdb;
  assign mem_MPORT_219_mask = 1'h1;
  assign mem_MPORT_219_en = reset;
  assign mem_MPORT_220_data = 32'h0;
  assign mem_MPORT_220_addr = 9'hdc;
  assign mem_MPORT_220_mask = 1'h1;
  assign mem_MPORT_220_en = reset;
  assign mem_MPORT_221_data = 32'h0;
  assign mem_MPORT_221_addr = 9'hdd;
  assign mem_MPORT_221_mask = 1'h1;
  assign mem_MPORT_221_en = reset;
  assign mem_MPORT_222_data = 32'h0;
  assign mem_MPORT_222_addr = 9'hde;
  assign mem_MPORT_222_mask = 1'h1;
  assign mem_MPORT_222_en = reset;
  assign mem_MPORT_223_data = 32'h0;
  assign mem_MPORT_223_addr = 9'hdf;
  assign mem_MPORT_223_mask = 1'h1;
  assign mem_MPORT_223_en = reset;
  assign mem_MPORT_224_data = 32'h0;
  assign mem_MPORT_224_addr = 9'he0;
  assign mem_MPORT_224_mask = 1'h1;
  assign mem_MPORT_224_en = reset;
  assign mem_MPORT_225_data = 32'h0;
  assign mem_MPORT_225_addr = 9'he1;
  assign mem_MPORT_225_mask = 1'h1;
  assign mem_MPORT_225_en = reset;
  assign mem_MPORT_226_data = 32'h0;
  assign mem_MPORT_226_addr = 9'he2;
  assign mem_MPORT_226_mask = 1'h1;
  assign mem_MPORT_226_en = reset;
  assign mem_MPORT_227_data = 32'h0;
  assign mem_MPORT_227_addr = 9'he3;
  assign mem_MPORT_227_mask = 1'h1;
  assign mem_MPORT_227_en = reset;
  assign mem_MPORT_228_data = 32'h0;
  assign mem_MPORT_228_addr = 9'he4;
  assign mem_MPORT_228_mask = 1'h1;
  assign mem_MPORT_228_en = reset;
  assign mem_MPORT_229_data = 32'h0;
  assign mem_MPORT_229_addr = 9'he5;
  assign mem_MPORT_229_mask = 1'h1;
  assign mem_MPORT_229_en = reset;
  assign mem_MPORT_230_data = 32'h0;
  assign mem_MPORT_230_addr = 9'he6;
  assign mem_MPORT_230_mask = 1'h1;
  assign mem_MPORT_230_en = reset;
  assign mem_MPORT_231_data = 32'h0;
  assign mem_MPORT_231_addr = 9'he7;
  assign mem_MPORT_231_mask = 1'h1;
  assign mem_MPORT_231_en = reset;
  assign mem_MPORT_232_data = 32'h0;
  assign mem_MPORT_232_addr = 9'he8;
  assign mem_MPORT_232_mask = 1'h1;
  assign mem_MPORT_232_en = reset;
  assign mem_MPORT_233_data = 32'h0;
  assign mem_MPORT_233_addr = 9'he9;
  assign mem_MPORT_233_mask = 1'h1;
  assign mem_MPORT_233_en = reset;
  assign mem_MPORT_234_data = 32'h0;
  assign mem_MPORT_234_addr = 9'hea;
  assign mem_MPORT_234_mask = 1'h1;
  assign mem_MPORT_234_en = reset;
  assign mem_MPORT_235_data = 32'h0;
  assign mem_MPORT_235_addr = 9'heb;
  assign mem_MPORT_235_mask = 1'h1;
  assign mem_MPORT_235_en = reset;
  assign mem_MPORT_236_data = 32'h0;
  assign mem_MPORT_236_addr = 9'hec;
  assign mem_MPORT_236_mask = 1'h1;
  assign mem_MPORT_236_en = reset;
  assign mem_MPORT_237_data = 32'h0;
  assign mem_MPORT_237_addr = 9'hed;
  assign mem_MPORT_237_mask = 1'h1;
  assign mem_MPORT_237_en = reset;
  assign mem_MPORT_238_data = 32'h0;
  assign mem_MPORT_238_addr = 9'hee;
  assign mem_MPORT_238_mask = 1'h1;
  assign mem_MPORT_238_en = reset;
  assign mem_MPORT_239_data = 32'h0;
  assign mem_MPORT_239_addr = 9'hef;
  assign mem_MPORT_239_mask = 1'h1;
  assign mem_MPORT_239_en = reset;
  assign mem_MPORT_240_data = 32'h0;
  assign mem_MPORT_240_addr = 9'hf0;
  assign mem_MPORT_240_mask = 1'h1;
  assign mem_MPORT_240_en = reset;
  assign mem_MPORT_241_data = 32'h0;
  assign mem_MPORT_241_addr = 9'hf1;
  assign mem_MPORT_241_mask = 1'h1;
  assign mem_MPORT_241_en = reset;
  assign mem_MPORT_242_data = 32'h0;
  assign mem_MPORT_242_addr = 9'hf2;
  assign mem_MPORT_242_mask = 1'h1;
  assign mem_MPORT_242_en = reset;
  assign mem_MPORT_243_data = 32'h0;
  assign mem_MPORT_243_addr = 9'hf3;
  assign mem_MPORT_243_mask = 1'h1;
  assign mem_MPORT_243_en = reset;
  assign mem_MPORT_244_data = 32'h0;
  assign mem_MPORT_244_addr = 9'hf4;
  assign mem_MPORT_244_mask = 1'h1;
  assign mem_MPORT_244_en = reset;
  assign mem_MPORT_245_data = 32'h0;
  assign mem_MPORT_245_addr = 9'hf5;
  assign mem_MPORT_245_mask = 1'h1;
  assign mem_MPORT_245_en = reset;
  assign mem_MPORT_246_data = 32'h0;
  assign mem_MPORT_246_addr = 9'hf6;
  assign mem_MPORT_246_mask = 1'h1;
  assign mem_MPORT_246_en = reset;
  assign mem_MPORT_247_data = 32'h0;
  assign mem_MPORT_247_addr = 9'hf7;
  assign mem_MPORT_247_mask = 1'h1;
  assign mem_MPORT_247_en = reset;
  assign mem_MPORT_248_data = 32'h0;
  assign mem_MPORT_248_addr = 9'hf8;
  assign mem_MPORT_248_mask = 1'h1;
  assign mem_MPORT_248_en = reset;
  assign mem_MPORT_249_data = 32'h0;
  assign mem_MPORT_249_addr = 9'hf9;
  assign mem_MPORT_249_mask = 1'h1;
  assign mem_MPORT_249_en = reset;
  assign mem_MPORT_250_data = 32'h0;
  assign mem_MPORT_250_addr = 9'hfa;
  assign mem_MPORT_250_mask = 1'h1;
  assign mem_MPORT_250_en = reset;
  assign mem_MPORT_251_data = 32'h0;
  assign mem_MPORT_251_addr = 9'hfb;
  assign mem_MPORT_251_mask = 1'h1;
  assign mem_MPORT_251_en = reset;
  assign mem_MPORT_252_data = 32'h0;
  assign mem_MPORT_252_addr = 9'hfc;
  assign mem_MPORT_252_mask = 1'h1;
  assign mem_MPORT_252_en = reset;
  assign mem_MPORT_253_data = 32'h0;
  assign mem_MPORT_253_addr = 9'hfd;
  assign mem_MPORT_253_mask = 1'h1;
  assign mem_MPORT_253_en = reset;
  assign mem_MPORT_254_data = 32'h0;
  assign mem_MPORT_254_addr = 9'hfe;
  assign mem_MPORT_254_mask = 1'h1;
  assign mem_MPORT_254_en = reset;
  assign mem_MPORT_255_data = 32'h0;
  assign mem_MPORT_255_addr = 9'hff;
  assign mem_MPORT_255_mask = 1'h1;
  assign mem_MPORT_255_en = reset;
  assign mem_MPORT_256_data = 32'h0;
  assign mem_MPORT_256_addr = 9'h100;
  assign mem_MPORT_256_mask = 1'h1;
  assign mem_MPORT_256_en = reset;
  assign mem_MPORT_257_data = 32'h0;
  assign mem_MPORT_257_addr = 9'h101;
  assign mem_MPORT_257_mask = 1'h1;
  assign mem_MPORT_257_en = reset;
  assign mem_MPORT_258_data = 32'h0;
  assign mem_MPORT_258_addr = 9'h102;
  assign mem_MPORT_258_mask = 1'h1;
  assign mem_MPORT_258_en = reset;
  assign mem_MPORT_259_data = 32'h0;
  assign mem_MPORT_259_addr = 9'h103;
  assign mem_MPORT_259_mask = 1'h1;
  assign mem_MPORT_259_en = reset;
  assign mem_MPORT_260_data = 32'h0;
  assign mem_MPORT_260_addr = 9'h104;
  assign mem_MPORT_260_mask = 1'h1;
  assign mem_MPORT_260_en = reset;
  assign mem_MPORT_261_data = 32'h0;
  assign mem_MPORT_261_addr = 9'h105;
  assign mem_MPORT_261_mask = 1'h1;
  assign mem_MPORT_261_en = reset;
  assign mem_MPORT_262_data = 32'h0;
  assign mem_MPORT_262_addr = 9'h106;
  assign mem_MPORT_262_mask = 1'h1;
  assign mem_MPORT_262_en = reset;
  assign mem_MPORT_263_data = 32'h0;
  assign mem_MPORT_263_addr = 9'h107;
  assign mem_MPORT_263_mask = 1'h1;
  assign mem_MPORT_263_en = reset;
  assign mem_MPORT_264_data = 32'h0;
  assign mem_MPORT_264_addr = 9'h108;
  assign mem_MPORT_264_mask = 1'h1;
  assign mem_MPORT_264_en = reset;
  assign mem_MPORT_265_data = 32'h0;
  assign mem_MPORT_265_addr = 9'h109;
  assign mem_MPORT_265_mask = 1'h1;
  assign mem_MPORT_265_en = reset;
  assign mem_MPORT_266_data = 32'h0;
  assign mem_MPORT_266_addr = 9'h10a;
  assign mem_MPORT_266_mask = 1'h1;
  assign mem_MPORT_266_en = reset;
  assign mem_MPORT_267_data = 32'h0;
  assign mem_MPORT_267_addr = 9'h10b;
  assign mem_MPORT_267_mask = 1'h1;
  assign mem_MPORT_267_en = reset;
  assign mem_MPORT_268_data = 32'h0;
  assign mem_MPORT_268_addr = 9'h10c;
  assign mem_MPORT_268_mask = 1'h1;
  assign mem_MPORT_268_en = reset;
  assign mem_MPORT_269_data = 32'h0;
  assign mem_MPORT_269_addr = 9'h10d;
  assign mem_MPORT_269_mask = 1'h1;
  assign mem_MPORT_269_en = reset;
  assign mem_MPORT_270_data = 32'h0;
  assign mem_MPORT_270_addr = 9'h10e;
  assign mem_MPORT_270_mask = 1'h1;
  assign mem_MPORT_270_en = reset;
  assign mem_MPORT_271_data = 32'h0;
  assign mem_MPORT_271_addr = 9'h10f;
  assign mem_MPORT_271_mask = 1'h1;
  assign mem_MPORT_271_en = reset;
  assign mem_MPORT_272_data = 32'h0;
  assign mem_MPORT_272_addr = 9'h110;
  assign mem_MPORT_272_mask = 1'h1;
  assign mem_MPORT_272_en = reset;
  assign mem_MPORT_273_data = 32'h0;
  assign mem_MPORT_273_addr = 9'h111;
  assign mem_MPORT_273_mask = 1'h1;
  assign mem_MPORT_273_en = reset;
  assign mem_MPORT_274_data = 32'h0;
  assign mem_MPORT_274_addr = 9'h112;
  assign mem_MPORT_274_mask = 1'h1;
  assign mem_MPORT_274_en = reset;
  assign mem_MPORT_275_data = 32'h0;
  assign mem_MPORT_275_addr = 9'h113;
  assign mem_MPORT_275_mask = 1'h1;
  assign mem_MPORT_275_en = reset;
  assign mem_MPORT_276_data = 32'h0;
  assign mem_MPORT_276_addr = 9'h114;
  assign mem_MPORT_276_mask = 1'h1;
  assign mem_MPORT_276_en = reset;
  assign mem_MPORT_277_data = 32'h0;
  assign mem_MPORT_277_addr = 9'h115;
  assign mem_MPORT_277_mask = 1'h1;
  assign mem_MPORT_277_en = reset;
  assign mem_MPORT_278_data = 32'h0;
  assign mem_MPORT_278_addr = 9'h116;
  assign mem_MPORT_278_mask = 1'h1;
  assign mem_MPORT_278_en = reset;
  assign mem_MPORT_279_data = 32'h0;
  assign mem_MPORT_279_addr = 9'h117;
  assign mem_MPORT_279_mask = 1'h1;
  assign mem_MPORT_279_en = reset;
  assign mem_MPORT_280_data = 32'h0;
  assign mem_MPORT_280_addr = 9'h118;
  assign mem_MPORT_280_mask = 1'h1;
  assign mem_MPORT_280_en = reset;
  assign mem_MPORT_281_data = 32'h0;
  assign mem_MPORT_281_addr = 9'h119;
  assign mem_MPORT_281_mask = 1'h1;
  assign mem_MPORT_281_en = reset;
  assign mem_MPORT_282_data = 32'h0;
  assign mem_MPORT_282_addr = 9'h11a;
  assign mem_MPORT_282_mask = 1'h1;
  assign mem_MPORT_282_en = reset;
  assign mem_MPORT_283_data = 32'h0;
  assign mem_MPORT_283_addr = 9'h11b;
  assign mem_MPORT_283_mask = 1'h1;
  assign mem_MPORT_283_en = reset;
  assign mem_MPORT_284_data = 32'h0;
  assign mem_MPORT_284_addr = 9'h11c;
  assign mem_MPORT_284_mask = 1'h1;
  assign mem_MPORT_284_en = reset;
  assign mem_MPORT_285_data = 32'h0;
  assign mem_MPORT_285_addr = 9'h11d;
  assign mem_MPORT_285_mask = 1'h1;
  assign mem_MPORT_285_en = reset;
  assign mem_MPORT_286_data = 32'h0;
  assign mem_MPORT_286_addr = 9'h11e;
  assign mem_MPORT_286_mask = 1'h1;
  assign mem_MPORT_286_en = reset;
  assign mem_MPORT_287_data = 32'h0;
  assign mem_MPORT_287_addr = 9'h11f;
  assign mem_MPORT_287_mask = 1'h1;
  assign mem_MPORT_287_en = reset;
  assign mem_MPORT_288_data = 32'h0;
  assign mem_MPORT_288_addr = 9'h120;
  assign mem_MPORT_288_mask = 1'h1;
  assign mem_MPORT_288_en = reset;
  assign mem_MPORT_289_data = 32'h0;
  assign mem_MPORT_289_addr = 9'h121;
  assign mem_MPORT_289_mask = 1'h1;
  assign mem_MPORT_289_en = reset;
  assign mem_MPORT_290_data = 32'h0;
  assign mem_MPORT_290_addr = 9'h122;
  assign mem_MPORT_290_mask = 1'h1;
  assign mem_MPORT_290_en = reset;
  assign mem_MPORT_291_data = 32'h0;
  assign mem_MPORT_291_addr = 9'h123;
  assign mem_MPORT_291_mask = 1'h1;
  assign mem_MPORT_291_en = reset;
  assign mem_MPORT_292_data = 32'h0;
  assign mem_MPORT_292_addr = 9'h124;
  assign mem_MPORT_292_mask = 1'h1;
  assign mem_MPORT_292_en = reset;
  assign mem_MPORT_293_data = 32'h0;
  assign mem_MPORT_293_addr = 9'h125;
  assign mem_MPORT_293_mask = 1'h1;
  assign mem_MPORT_293_en = reset;
  assign mem_MPORT_294_data = 32'h0;
  assign mem_MPORT_294_addr = 9'h126;
  assign mem_MPORT_294_mask = 1'h1;
  assign mem_MPORT_294_en = reset;
  assign mem_MPORT_295_data = 32'h0;
  assign mem_MPORT_295_addr = 9'h127;
  assign mem_MPORT_295_mask = 1'h1;
  assign mem_MPORT_295_en = reset;
  assign mem_MPORT_296_data = 32'h0;
  assign mem_MPORT_296_addr = 9'h128;
  assign mem_MPORT_296_mask = 1'h1;
  assign mem_MPORT_296_en = reset;
  assign mem_MPORT_297_data = 32'h0;
  assign mem_MPORT_297_addr = 9'h129;
  assign mem_MPORT_297_mask = 1'h1;
  assign mem_MPORT_297_en = reset;
  assign mem_MPORT_298_data = 32'h0;
  assign mem_MPORT_298_addr = 9'h12a;
  assign mem_MPORT_298_mask = 1'h1;
  assign mem_MPORT_298_en = reset;
  assign mem_MPORT_299_data = 32'h0;
  assign mem_MPORT_299_addr = 9'h12b;
  assign mem_MPORT_299_mask = 1'h1;
  assign mem_MPORT_299_en = reset;
  assign mem_MPORT_300_data = 32'h0;
  assign mem_MPORT_300_addr = 9'h12c;
  assign mem_MPORT_300_mask = 1'h1;
  assign mem_MPORT_300_en = reset;
  assign mem_MPORT_301_data = 32'h0;
  assign mem_MPORT_301_addr = 9'h12d;
  assign mem_MPORT_301_mask = 1'h1;
  assign mem_MPORT_301_en = reset;
  assign mem_MPORT_302_data = 32'h0;
  assign mem_MPORT_302_addr = 9'h12e;
  assign mem_MPORT_302_mask = 1'h1;
  assign mem_MPORT_302_en = reset;
  assign mem_MPORT_303_data = 32'h0;
  assign mem_MPORT_303_addr = 9'h12f;
  assign mem_MPORT_303_mask = 1'h1;
  assign mem_MPORT_303_en = reset;
  assign mem_MPORT_304_data = 32'h0;
  assign mem_MPORT_304_addr = 9'h130;
  assign mem_MPORT_304_mask = 1'h1;
  assign mem_MPORT_304_en = reset;
  assign mem_MPORT_305_data = 32'h0;
  assign mem_MPORT_305_addr = 9'h131;
  assign mem_MPORT_305_mask = 1'h1;
  assign mem_MPORT_305_en = reset;
  assign mem_MPORT_306_data = 32'h0;
  assign mem_MPORT_306_addr = 9'h132;
  assign mem_MPORT_306_mask = 1'h1;
  assign mem_MPORT_306_en = reset;
  assign mem_MPORT_307_data = 32'h0;
  assign mem_MPORT_307_addr = 9'h133;
  assign mem_MPORT_307_mask = 1'h1;
  assign mem_MPORT_307_en = reset;
  assign mem_MPORT_308_data = 32'h0;
  assign mem_MPORT_308_addr = 9'h134;
  assign mem_MPORT_308_mask = 1'h1;
  assign mem_MPORT_308_en = reset;
  assign mem_MPORT_309_data = 32'h0;
  assign mem_MPORT_309_addr = 9'h135;
  assign mem_MPORT_309_mask = 1'h1;
  assign mem_MPORT_309_en = reset;
  assign mem_MPORT_310_data = 32'h0;
  assign mem_MPORT_310_addr = 9'h136;
  assign mem_MPORT_310_mask = 1'h1;
  assign mem_MPORT_310_en = reset;
  assign mem_MPORT_311_data = 32'h0;
  assign mem_MPORT_311_addr = 9'h137;
  assign mem_MPORT_311_mask = 1'h1;
  assign mem_MPORT_311_en = reset;
  assign mem_MPORT_312_data = 32'h0;
  assign mem_MPORT_312_addr = 9'h138;
  assign mem_MPORT_312_mask = 1'h1;
  assign mem_MPORT_312_en = reset;
  assign mem_MPORT_313_data = 32'h0;
  assign mem_MPORT_313_addr = 9'h139;
  assign mem_MPORT_313_mask = 1'h1;
  assign mem_MPORT_313_en = reset;
  assign mem_MPORT_314_data = 32'h0;
  assign mem_MPORT_314_addr = 9'h13a;
  assign mem_MPORT_314_mask = 1'h1;
  assign mem_MPORT_314_en = reset;
  assign mem_MPORT_315_data = 32'h0;
  assign mem_MPORT_315_addr = 9'h13b;
  assign mem_MPORT_315_mask = 1'h1;
  assign mem_MPORT_315_en = reset;
  assign mem_MPORT_316_data = 32'h0;
  assign mem_MPORT_316_addr = 9'h13c;
  assign mem_MPORT_316_mask = 1'h1;
  assign mem_MPORT_316_en = reset;
  assign mem_MPORT_317_data = 32'h0;
  assign mem_MPORT_317_addr = 9'h13d;
  assign mem_MPORT_317_mask = 1'h1;
  assign mem_MPORT_317_en = reset;
  assign mem_MPORT_318_data = 32'h0;
  assign mem_MPORT_318_addr = 9'h13e;
  assign mem_MPORT_318_mask = 1'h1;
  assign mem_MPORT_318_en = reset;
  assign mem_MPORT_319_data = 32'h0;
  assign mem_MPORT_319_addr = 9'h13f;
  assign mem_MPORT_319_mask = 1'h1;
  assign mem_MPORT_319_en = reset;
  assign mem_MPORT_320_data = 32'h0;
  assign mem_MPORT_320_addr = 9'h140;
  assign mem_MPORT_320_mask = 1'h1;
  assign mem_MPORT_320_en = reset;
  assign mem_MPORT_321_data = 32'h0;
  assign mem_MPORT_321_addr = 9'h141;
  assign mem_MPORT_321_mask = 1'h1;
  assign mem_MPORT_321_en = reset;
  assign mem_MPORT_322_data = 32'h0;
  assign mem_MPORT_322_addr = 9'h142;
  assign mem_MPORT_322_mask = 1'h1;
  assign mem_MPORT_322_en = reset;
  assign mem_MPORT_323_data = 32'h0;
  assign mem_MPORT_323_addr = 9'h143;
  assign mem_MPORT_323_mask = 1'h1;
  assign mem_MPORT_323_en = reset;
  assign mem_MPORT_324_data = 32'h0;
  assign mem_MPORT_324_addr = 9'h144;
  assign mem_MPORT_324_mask = 1'h1;
  assign mem_MPORT_324_en = reset;
  assign mem_MPORT_325_data = 32'h0;
  assign mem_MPORT_325_addr = 9'h145;
  assign mem_MPORT_325_mask = 1'h1;
  assign mem_MPORT_325_en = reset;
  assign mem_MPORT_326_data = 32'h0;
  assign mem_MPORT_326_addr = 9'h146;
  assign mem_MPORT_326_mask = 1'h1;
  assign mem_MPORT_326_en = reset;
  assign mem_MPORT_327_data = 32'h0;
  assign mem_MPORT_327_addr = 9'h147;
  assign mem_MPORT_327_mask = 1'h1;
  assign mem_MPORT_327_en = reset;
  assign mem_MPORT_328_data = 32'h0;
  assign mem_MPORT_328_addr = 9'h148;
  assign mem_MPORT_328_mask = 1'h1;
  assign mem_MPORT_328_en = reset;
  assign mem_MPORT_329_data = 32'h0;
  assign mem_MPORT_329_addr = 9'h149;
  assign mem_MPORT_329_mask = 1'h1;
  assign mem_MPORT_329_en = reset;
  assign mem_MPORT_330_data = 32'h0;
  assign mem_MPORT_330_addr = 9'h14a;
  assign mem_MPORT_330_mask = 1'h1;
  assign mem_MPORT_330_en = reset;
  assign mem_MPORT_331_data = 32'h0;
  assign mem_MPORT_331_addr = 9'h14b;
  assign mem_MPORT_331_mask = 1'h1;
  assign mem_MPORT_331_en = reset;
  assign mem_MPORT_332_data = 32'h0;
  assign mem_MPORT_332_addr = 9'h14c;
  assign mem_MPORT_332_mask = 1'h1;
  assign mem_MPORT_332_en = reset;
  assign mem_MPORT_333_data = 32'h0;
  assign mem_MPORT_333_addr = 9'h14d;
  assign mem_MPORT_333_mask = 1'h1;
  assign mem_MPORT_333_en = reset;
  assign mem_MPORT_334_data = 32'h0;
  assign mem_MPORT_334_addr = 9'h14e;
  assign mem_MPORT_334_mask = 1'h1;
  assign mem_MPORT_334_en = reset;
  assign mem_MPORT_335_data = 32'h0;
  assign mem_MPORT_335_addr = 9'h14f;
  assign mem_MPORT_335_mask = 1'h1;
  assign mem_MPORT_335_en = reset;
  assign mem_MPORT_336_data = 32'h0;
  assign mem_MPORT_336_addr = 9'h150;
  assign mem_MPORT_336_mask = 1'h1;
  assign mem_MPORT_336_en = reset;
  assign mem_MPORT_337_data = 32'h0;
  assign mem_MPORT_337_addr = 9'h151;
  assign mem_MPORT_337_mask = 1'h1;
  assign mem_MPORT_337_en = reset;
  assign mem_MPORT_338_data = 32'h0;
  assign mem_MPORT_338_addr = 9'h152;
  assign mem_MPORT_338_mask = 1'h1;
  assign mem_MPORT_338_en = reset;
  assign mem_MPORT_339_data = 32'h0;
  assign mem_MPORT_339_addr = 9'h153;
  assign mem_MPORT_339_mask = 1'h1;
  assign mem_MPORT_339_en = reset;
  assign mem_MPORT_340_data = 32'h0;
  assign mem_MPORT_340_addr = 9'h154;
  assign mem_MPORT_340_mask = 1'h1;
  assign mem_MPORT_340_en = reset;
  assign mem_MPORT_341_data = 32'h0;
  assign mem_MPORT_341_addr = 9'h155;
  assign mem_MPORT_341_mask = 1'h1;
  assign mem_MPORT_341_en = reset;
  assign mem_MPORT_342_data = 32'h0;
  assign mem_MPORT_342_addr = 9'h156;
  assign mem_MPORT_342_mask = 1'h1;
  assign mem_MPORT_342_en = reset;
  assign mem_MPORT_343_data = 32'h0;
  assign mem_MPORT_343_addr = 9'h157;
  assign mem_MPORT_343_mask = 1'h1;
  assign mem_MPORT_343_en = reset;
  assign mem_MPORT_344_data = 32'h0;
  assign mem_MPORT_344_addr = 9'h158;
  assign mem_MPORT_344_mask = 1'h1;
  assign mem_MPORT_344_en = reset;
  assign mem_MPORT_345_data = 32'h0;
  assign mem_MPORT_345_addr = 9'h159;
  assign mem_MPORT_345_mask = 1'h1;
  assign mem_MPORT_345_en = reset;
  assign mem_MPORT_346_data = 32'h0;
  assign mem_MPORT_346_addr = 9'h15a;
  assign mem_MPORT_346_mask = 1'h1;
  assign mem_MPORT_346_en = reset;
  assign mem_MPORT_347_data = 32'h0;
  assign mem_MPORT_347_addr = 9'h15b;
  assign mem_MPORT_347_mask = 1'h1;
  assign mem_MPORT_347_en = reset;
  assign mem_MPORT_348_data = 32'h0;
  assign mem_MPORT_348_addr = 9'h15c;
  assign mem_MPORT_348_mask = 1'h1;
  assign mem_MPORT_348_en = reset;
  assign mem_MPORT_349_data = 32'h0;
  assign mem_MPORT_349_addr = 9'h15d;
  assign mem_MPORT_349_mask = 1'h1;
  assign mem_MPORT_349_en = reset;
  assign mem_MPORT_350_data = 32'h0;
  assign mem_MPORT_350_addr = 9'h15e;
  assign mem_MPORT_350_mask = 1'h1;
  assign mem_MPORT_350_en = reset;
  assign mem_MPORT_351_data = 32'h0;
  assign mem_MPORT_351_addr = 9'h15f;
  assign mem_MPORT_351_mask = 1'h1;
  assign mem_MPORT_351_en = reset;
  assign mem_MPORT_352_data = 32'h0;
  assign mem_MPORT_352_addr = 9'h160;
  assign mem_MPORT_352_mask = 1'h1;
  assign mem_MPORT_352_en = reset;
  assign mem_MPORT_353_data = 32'h0;
  assign mem_MPORT_353_addr = 9'h161;
  assign mem_MPORT_353_mask = 1'h1;
  assign mem_MPORT_353_en = reset;
  assign mem_MPORT_354_data = 32'h0;
  assign mem_MPORT_354_addr = 9'h162;
  assign mem_MPORT_354_mask = 1'h1;
  assign mem_MPORT_354_en = reset;
  assign mem_MPORT_355_data = 32'h0;
  assign mem_MPORT_355_addr = 9'h163;
  assign mem_MPORT_355_mask = 1'h1;
  assign mem_MPORT_355_en = reset;
  assign mem_MPORT_356_data = 32'h0;
  assign mem_MPORT_356_addr = 9'h164;
  assign mem_MPORT_356_mask = 1'h1;
  assign mem_MPORT_356_en = reset;
  assign mem_MPORT_357_data = 32'h0;
  assign mem_MPORT_357_addr = 9'h165;
  assign mem_MPORT_357_mask = 1'h1;
  assign mem_MPORT_357_en = reset;
  assign mem_MPORT_358_data = 32'h0;
  assign mem_MPORT_358_addr = 9'h166;
  assign mem_MPORT_358_mask = 1'h1;
  assign mem_MPORT_358_en = reset;
  assign mem_MPORT_359_data = 32'h0;
  assign mem_MPORT_359_addr = 9'h167;
  assign mem_MPORT_359_mask = 1'h1;
  assign mem_MPORT_359_en = reset;
  assign mem_MPORT_360_data = 32'h0;
  assign mem_MPORT_360_addr = 9'h168;
  assign mem_MPORT_360_mask = 1'h1;
  assign mem_MPORT_360_en = reset;
  assign mem_MPORT_361_data = 32'h0;
  assign mem_MPORT_361_addr = 9'h169;
  assign mem_MPORT_361_mask = 1'h1;
  assign mem_MPORT_361_en = reset;
  assign mem_MPORT_362_data = 32'h0;
  assign mem_MPORT_362_addr = 9'h16a;
  assign mem_MPORT_362_mask = 1'h1;
  assign mem_MPORT_362_en = reset;
  assign mem_MPORT_363_data = 32'h0;
  assign mem_MPORT_363_addr = 9'h16b;
  assign mem_MPORT_363_mask = 1'h1;
  assign mem_MPORT_363_en = reset;
  assign mem_MPORT_364_data = 32'h0;
  assign mem_MPORT_364_addr = 9'h16c;
  assign mem_MPORT_364_mask = 1'h1;
  assign mem_MPORT_364_en = reset;
  assign mem_MPORT_365_data = 32'h0;
  assign mem_MPORT_365_addr = 9'h16d;
  assign mem_MPORT_365_mask = 1'h1;
  assign mem_MPORT_365_en = reset;
  assign mem_MPORT_366_data = 32'h0;
  assign mem_MPORT_366_addr = 9'h16e;
  assign mem_MPORT_366_mask = 1'h1;
  assign mem_MPORT_366_en = reset;
  assign mem_MPORT_367_data = 32'h0;
  assign mem_MPORT_367_addr = 9'h16f;
  assign mem_MPORT_367_mask = 1'h1;
  assign mem_MPORT_367_en = reset;
  assign mem_MPORT_368_data = 32'h0;
  assign mem_MPORT_368_addr = 9'h170;
  assign mem_MPORT_368_mask = 1'h1;
  assign mem_MPORT_368_en = reset;
  assign mem_MPORT_369_data = 32'h0;
  assign mem_MPORT_369_addr = 9'h171;
  assign mem_MPORT_369_mask = 1'h1;
  assign mem_MPORT_369_en = reset;
  assign mem_MPORT_370_data = 32'h0;
  assign mem_MPORT_370_addr = 9'h172;
  assign mem_MPORT_370_mask = 1'h1;
  assign mem_MPORT_370_en = reset;
  assign mem_MPORT_371_data = 32'h0;
  assign mem_MPORT_371_addr = 9'h173;
  assign mem_MPORT_371_mask = 1'h1;
  assign mem_MPORT_371_en = reset;
  assign mem_MPORT_372_data = 32'h0;
  assign mem_MPORT_372_addr = 9'h174;
  assign mem_MPORT_372_mask = 1'h1;
  assign mem_MPORT_372_en = reset;
  assign mem_MPORT_373_data = 32'h0;
  assign mem_MPORT_373_addr = 9'h175;
  assign mem_MPORT_373_mask = 1'h1;
  assign mem_MPORT_373_en = reset;
  assign mem_MPORT_374_data = 32'h0;
  assign mem_MPORT_374_addr = 9'h176;
  assign mem_MPORT_374_mask = 1'h1;
  assign mem_MPORT_374_en = reset;
  assign mem_MPORT_375_data = 32'h0;
  assign mem_MPORT_375_addr = 9'h177;
  assign mem_MPORT_375_mask = 1'h1;
  assign mem_MPORT_375_en = reset;
  assign mem_MPORT_376_data = 32'h0;
  assign mem_MPORT_376_addr = 9'h178;
  assign mem_MPORT_376_mask = 1'h1;
  assign mem_MPORT_376_en = reset;
  assign mem_MPORT_377_data = 32'h0;
  assign mem_MPORT_377_addr = 9'h179;
  assign mem_MPORT_377_mask = 1'h1;
  assign mem_MPORT_377_en = reset;
  assign mem_MPORT_378_data = 32'h0;
  assign mem_MPORT_378_addr = 9'h17a;
  assign mem_MPORT_378_mask = 1'h1;
  assign mem_MPORT_378_en = reset;
  assign mem_MPORT_379_data = 32'h0;
  assign mem_MPORT_379_addr = 9'h17b;
  assign mem_MPORT_379_mask = 1'h1;
  assign mem_MPORT_379_en = reset;
  assign mem_MPORT_380_data = 32'h0;
  assign mem_MPORT_380_addr = 9'h17c;
  assign mem_MPORT_380_mask = 1'h1;
  assign mem_MPORT_380_en = reset;
  assign mem_MPORT_381_data = 32'h0;
  assign mem_MPORT_381_addr = 9'h17d;
  assign mem_MPORT_381_mask = 1'h1;
  assign mem_MPORT_381_en = reset;
  assign mem_MPORT_382_data = 32'h0;
  assign mem_MPORT_382_addr = 9'h17e;
  assign mem_MPORT_382_mask = 1'h1;
  assign mem_MPORT_382_en = reset;
  assign mem_MPORT_383_data = 32'h0;
  assign mem_MPORT_383_addr = 9'h17f;
  assign mem_MPORT_383_mask = 1'h1;
  assign mem_MPORT_383_en = reset;
  assign mem_MPORT_384_data = 32'h0;
  assign mem_MPORT_384_addr = 9'h180;
  assign mem_MPORT_384_mask = 1'h1;
  assign mem_MPORT_384_en = reset;
  assign mem_MPORT_385_data = 32'h0;
  assign mem_MPORT_385_addr = 9'h181;
  assign mem_MPORT_385_mask = 1'h1;
  assign mem_MPORT_385_en = reset;
  assign mem_MPORT_386_data = 32'h0;
  assign mem_MPORT_386_addr = 9'h182;
  assign mem_MPORT_386_mask = 1'h1;
  assign mem_MPORT_386_en = reset;
  assign mem_MPORT_387_data = 32'h0;
  assign mem_MPORT_387_addr = 9'h183;
  assign mem_MPORT_387_mask = 1'h1;
  assign mem_MPORT_387_en = reset;
  assign mem_MPORT_388_data = 32'h0;
  assign mem_MPORT_388_addr = 9'h184;
  assign mem_MPORT_388_mask = 1'h1;
  assign mem_MPORT_388_en = reset;
  assign mem_MPORT_389_data = 32'h0;
  assign mem_MPORT_389_addr = 9'h185;
  assign mem_MPORT_389_mask = 1'h1;
  assign mem_MPORT_389_en = reset;
  assign mem_MPORT_390_data = 32'h0;
  assign mem_MPORT_390_addr = 9'h186;
  assign mem_MPORT_390_mask = 1'h1;
  assign mem_MPORT_390_en = reset;
  assign mem_MPORT_391_data = 32'h0;
  assign mem_MPORT_391_addr = 9'h187;
  assign mem_MPORT_391_mask = 1'h1;
  assign mem_MPORT_391_en = reset;
  assign mem_MPORT_392_data = 32'h0;
  assign mem_MPORT_392_addr = 9'h188;
  assign mem_MPORT_392_mask = 1'h1;
  assign mem_MPORT_392_en = reset;
  assign mem_MPORT_393_data = 32'h0;
  assign mem_MPORT_393_addr = 9'h189;
  assign mem_MPORT_393_mask = 1'h1;
  assign mem_MPORT_393_en = reset;
  assign mem_MPORT_394_data = 32'h0;
  assign mem_MPORT_394_addr = 9'h18a;
  assign mem_MPORT_394_mask = 1'h1;
  assign mem_MPORT_394_en = reset;
  assign mem_MPORT_395_data = 32'h0;
  assign mem_MPORT_395_addr = 9'h18b;
  assign mem_MPORT_395_mask = 1'h1;
  assign mem_MPORT_395_en = reset;
  assign mem_MPORT_396_data = 32'h0;
  assign mem_MPORT_396_addr = 9'h18c;
  assign mem_MPORT_396_mask = 1'h1;
  assign mem_MPORT_396_en = reset;
  assign mem_MPORT_397_data = 32'h0;
  assign mem_MPORT_397_addr = 9'h18d;
  assign mem_MPORT_397_mask = 1'h1;
  assign mem_MPORT_397_en = reset;
  assign mem_MPORT_398_data = 32'h0;
  assign mem_MPORT_398_addr = 9'h18e;
  assign mem_MPORT_398_mask = 1'h1;
  assign mem_MPORT_398_en = reset;
  assign mem_MPORT_399_data = 32'h0;
  assign mem_MPORT_399_addr = 9'h18f;
  assign mem_MPORT_399_mask = 1'h1;
  assign mem_MPORT_399_en = reset;
  assign mem_MPORT_400_data = 32'h0;
  assign mem_MPORT_400_addr = 9'h190;
  assign mem_MPORT_400_mask = 1'h1;
  assign mem_MPORT_400_en = reset;
  assign mem_MPORT_401_data = 32'h0;
  assign mem_MPORT_401_addr = 9'h191;
  assign mem_MPORT_401_mask = 1'h1;
  assign mem_MPORT_401_en = reset;
  assign mem_MPORT_402_data = 32'h0;
  assign mem_MPORT_402_addr = 9'h192;
  assign mem_MPORT_402_mask = 1'h1;
  assign mem_MPORT_402_en = reset;
  assign mem_MPORT_403_data = 32'h0;
  assign mem_MPORT_403_addr = 9'h193;
  assign mem_MPORT_403_mask = 1'h1;
  assign mem_MPORT_403_en = reset;
  assign mem_MPORT_404_data = 32'h0;
  assign mem_MPORT_404_addr = 9'h194;
  assign mem_MPORT_404_mask = 1'h1;
  assign mem_MPORT_404_en = reset;
  assign mem_MPORT_405_data = 32'h0;
  assign mem_MPORT_405_addr = 9'h195;
  assign mem_MPORT_405_mask = 1'h1;
  assign mem_MPORT_405_en = reset;
  assign mem_MPORT_406_data = 32'h0;
  assign mem_MPORT_406_addr = 9'h196;
  assign mem_MPORT_406_mask = 1'h1;
  assign mem_MPORT_406_en = reset;
  assign mem_MPORT_407_data = 32'h0;
  assign mem_MPORT_407_addr = 9'h197;
  assign mem_MPORT_407_mask = 1'h1;
  assign mem_MPORT_407_en = reset;
  assign mem_MPORT_408_data = 32'h0;
  assign mem_MPORT_408_addr = 9'h198;
  assign mem_MPORT_408_mask = 1'h1;
  assign mem_MPORT_408_en = reset;
  assign mem_MPORT_409_data = 32'h0;
  assign mem_MPORT_409_addr = 9'h199;
  assign mem_MPORT_409_mask = 1'h1;
  assign mem_MPORT_409_en = reset;
  assign mem_MPORT_410_data = 32'h0;
  assign mem_MPORT_410_addr = 9'h19a;
  assign mem_MPORT_410_mask = 1'h1;
  assign mem_MPORT_410_en = reset;
  assign mem_MPORT_411_data = 32'h0;
  assign mem_MPORT_411_addr = 9'h19b;
  assign mem_MPORT_411_mask = 1'h1;
  assign mem_MPORT_411_en = reset;
  assign mem_MPORT_412_data = 32'h0;
  assign mem_MPORT_412_addr = 9'h19c;
  assign mem_MPORT_412_mask = 1'h1;
  assign mem_MPORT_412_en = reset;
  assign mem_MPORT_413_data = 32'h0;
  assign mem_MPORT_413_addr = 9'h19d;
  assign mem_MPORT_413_mask = 1'h1;
  assign mem_MPORT_413_en = reset;
  assign mem_MPORT_414_data = 32'h0;
  assign mem_MPORT_414_addr = 9'h19e;
  assign mem_MPORT_414_mask = 1'h1;
  assign mem_MPORT_414_en = reset;
  assign mem_MPORT_415_data = 32'h0;
  assign mem_MPORT_415_addr = 9'h19f;
  assign mem_MPORT_415_mask = 1'h1;
  assign mem_MPORT_415_en = reset;
  assign mem_MPORT_416_data = 32'h0;
  assign mem_MPORT_416_addr = 9'h1a0;
  assign mem_MPORT_416_mask = 1'h1;
  assign mem_MPORT_416_en = reset;
  assign mem_MPORT_417_data = 32'h0;
  assign mem_MPORT_417_addr = 9'h1a1;
  assign mem_MPORT_417_mask = 1'h1;
  assign mem_MPORT_417_en = reset;
  assign mem_MPORT_418_data = 32'h0;
  assign mem_MPORT_418_addr = 9'h1a2;
  assign mem_MPORT_418_mask = 1'h1;
  assign mem_MPORT_418_en = reset;
  assign mem_MPORT_419_data = 32'h0;
  assign mem_MPORT_419_addr = 9'h1a3;
  assign mem_MPORT_419_mask = 1'h1;
  assign mem_MPORT_419_en = reset;
  assign mem_MPORT_420_data = 32'h0;
  assign mem_MPORT_420_addr = 9'h1a4;
  assign mem_MPORT_420_mask = 1'h1;
  assign mem_MPORT_420_en = reset;
  assign mem_MPORT_421_data = 32'h0;
  assign mem_MPORT_421_addr = 9'h1a5;
  assign mem_MPORT_421_mask = 1'h1;
  assign mem_MPORT_421_en = reset;
  assign mem_MPORT_422_data = 32'h0;
  assign mem_MPORT_422_addr = 9'h1a6;
  assign mem_MPORT_422_mask = 1'h1;
  assign mem_MPORT_422_en = reset;
  assign mem_MPORT_423_data = 32'h0;
  assign mem_MPORT_423_addr = 9'h1a7;
  assign mem_MPORT_423_mask = 1'h1;
  assign mem_MPORT_423_en = reset;
  assign mem_MPORT_424_data = 32'h0;
  assign mem_MPORT_424_addr = 9'h1a8;
  assign mem_MPORT_424_mask = 1'h1;
  assign mem_MPORT_424_en = reset;
  assign mem_MPORT_425_data = 32'h0;
  assign mem_MPORT_425_addr = 9'h1a9;
  assign mem_MPORT_425_mask = 1'h1;
  assign mem_MPORT_425_en = reset;
  assign mem_MPORT_426_data = 32'h0;
  assign mem_MPORT_426_addr = 9'h1aa;
  assign mem_MPORT_426_mask = 1'h1;
  assign mem_MPORT_426_en = reset;
  assign mem_MPORT_427_data = 32'h0;
  assign mem_MPORT_427_addr = 9'h1ab;
  assign mem_MPORT_427_mask = 1'h1;
  assign mem_MPORT_427_en = reset;
  assign mem_MPORT_428_data = 32'h0;
  assign mem_MPORT_428_addr = 9'h1ac;
  assign mem_MPORT_428_mask = 1'h1;
  assign mem_MPORT_428_en = reset;
  assign mem_MPORT_429_data = 32'h0;
  assign mem_MPORT_429_addr = 9'h1ad;
  assign mem_MPORT_429_mask = 1'h1;
  assign mem_MPORT_429_en = reset;
  assign mem_MPORT_430_data = 32'h0;
  assign mem_MPORT_430_addr = 9'h1ae;
  assign mem_MPORT_430_mask = 1'h1;
  assign mem_MPORT_430_en = reset;
  assign mem_MPORT_431_data = 32'h0;
  assign mem_MPORT_431_addr = 9'h1af;
  assign mem_MPORT_431_mask = 1'h1;
  assign mem_MPORT_431_en = reset;
  assign mem_MPORT_432_data = 32'h0;
  assign mem_MPORT_432_addr = 9'h1b0;
  assign mem_MPORT_432_mask = 1'h1;
  assign mem_MPORT_432_en = reset;
  assign mem_MPORT_433_data = 32'h0;
  assign mem_MPORT_433_addr = 9'h1b1;
  assign mem_MPORT_433_mask = 1'h1;
  assign mem_MPORT_433_en = reset;
  assign mem_MPORT_434_data = 32'h0;
  assign mem_MPORT_434_addr = 9'h1b2;
  assign mem_MPORT_434_mask = 1'h1;
  assign mem_MPORT_434_en = reset;
  assign mem_MPORT_435_data = 32'h0;
  assign mem_MPORT_435_addr = 9'h1b3;
  assign mem_MPORT_435_mask = 1'h1;
  assign mem_MPORT_435_en = reset;
  assign mem_MPORT_436_data = 32'h0;
  assign mem_MPORT_436_addr = 9'h1b4;
  assign mem_MPORT_436_mask = 1'h1;
  assign mem_MPORT_436_en = reset;
  assign mem_MPORT_437_data = 32'h0;
  assign mem_MPORT_437_addr = 9'h1b5;
  assign mem_MPORT_437_mask = 1'h1;
  assign mem_MPORT_437_en = reset;
  assign mem_MPORT_438_data = 32'h0;
  assign mem_MPORT_438_addr = 9'h1b6;
  assign mem_MPORT_438_mask = 1'h1;
  assign mem_MPORT_438_en = reset;
  assign mem_MPORT_439_data = 32'h0;
  assign mem_MPORT_439_addr = 9'h1b7;
  assign mem_MPORT_439_mask = 1'h1;
  assign mem_MPORT_439_en = reset;
  assign mem_MPORT_440_data = 32'h0;
  assign mem_MPORT_440_addr = 9'h1b8;
  assign mem_MPORT_440_mask = 1'h1;
  assign mem_MPORT_440_en = reset;
  assign mem_MPORT_441_data = 32'h0;
  assign mem_MPORT_441_addr = 9'h1b9;
  assign mem_MPORT_441_mask = 1'h1;
  assign mem_MPORT_441_en = reset;
  assign mem_MPORT_442_data = 32'h0;
  assign mem_MPORT_442_addr = 9'h1ba;
  assign mem_MPORT_442_mask = 1'h1;
  assign mem_MPORT_442_en = reset;
  assign mem_MPORT_443_data = 32'h0;
  assign mem_MPORT_443_addr = 9'h1bb;
  assign mem_MPORT_443_mask = 1'h1;
  assign mem_MPORT_443_en = reset;
  assign mem_MPORT_444_data = 32'h0;
  assign mem_MPORT_444_addr = 9'h1bc;
  assign mem_MPORT_444_mask = 1'h1;
  assign mem_MPORT_444_en = reset;
  assign mem_MPORT_445_data = 32'h0;
  assign mem_MPORT_445_addr = 9'h1bd;
  assign mem_MPORT_445_mask = 1'h1;
  assign mem_MPORT_445_en = reset;
  assign mem_MPORT_446_data = 32'h0;
  assign mem_MPORT_446_addr = 9'h1be;
  assign mem_MPORT_446_mask = 1'h1;
  assign mem_MPORT_446_en = reset;
  assign mem_MPORT_447_data = 32'h0;
  assign mem_MPORT_447_addr = 9'h1bf;
  assign mem_MPORT_447_mask = 1'h1;
  assign mem_MPORT_447_en = reset;
  assign mem_MPORT_448_data = 32'h0;
  assign mem_MPORT_448_addr = 9'h1c0;
  assign mem_MPORT_448_mask = 1'h1;
  assign mem_MPORT_448_en = reset;
  assign mem_MPORT_449_data = 32'h0;
  assign mem_MPORT_449_addr = 9'h1c1;
  assign mem_MPORT_449_mask = 1'h1;
  assign mem_MPORT_449_en = reset;
  assign mem_MPORT_450_data = 32'h0;
  assign mem_MPORT_450_addr = 9'h1c2;
  assign mem_MPORT_450_mask = 1'h1;
  assign mem_MPORT_450_en = reset;
  assign mem_MPORT_451_data = 32'h0;
  assign mem_MPORT_451_addr = 9'h1c3;
  assign mem_MPORT_451_mask = 1'h1;
  assign mem_MPORT_451_en = reset;
  assign mem_MPORT_452_data = 32'h0;
  assign mem_MPORT_452_addr = 9'h1c4;
  assign mem_MPORT_452_mask = 1'h1;
  assign mem_MPORT_452_en = reset;
  assign mem_MPORT_453_data = 32'h0;
  assign mem_MPORT_453_addr = 9'h1c5;
  assign mem_MPORT_453_mask = 1'h1;
  assign mem_MPORT_453_en = reset;
  assign mem_MPORT_454_data = 32'h0;
  assign mem_MPORT_454_addr = 9'h1c6;
  assign mem_MPORT_454_mask = 1'h1;
  assign mem_MPORT_454_en = reset;
  assign mem_MPORT_455_data = 32'h0;
  assign mem_MPORT_455_addr = 9'h1c7;
  assign mem_MPORT_455_mask = 1'h1;
  assign mem_MPORT_455_en = reset;
  assign mem_MPORT_456_data = 32'h0;
  assign mem_MPORT_456_addr = 9'h1c8;
  assign mem_MPORT_456_mask = 1'h1;
  assign mem_MPORT_456_en = reset;
  assign mem_MPORT_457_data = 32'h0;
  assign mem_MPORT_457_addr = 9'h1c9;
  assign mem_MPORT_457_mask = 1'h1;
  assign mem_MPORT_457_en = reset;
  assign mem_MPORT_458_data = 32'h0;
  assign mem_MPORT_458_addr = 9'h1ca;
  assign mem_MPORT_458_mask = 1'h1;
  assign mem_MPORT_458_en = reset;
  assign mem_MPORT_459_data = 32'h0;
  assign mem_MPORT_459_addr = 9'h1cb;
  assign mem_MPORT_459_mask = 1'h1;
  assign mem_MPORT_459_en = reset;
  assign mem_MPORT_460_data = 32'h0;
  assign mem_MPORT_460_addr = 9'h1cc;
  assign mem_MPORT_460_mask = 1'h1;
  assign mem_MPORT_460_en = reset;
  assign mem_MPORT_461_data = 32'h0;
  assign mem_MPORT_461_addr = 9'h1cd;
  assign mem_MPORT_461_mask = 1'h1;
  assign mem_MPORT_461_en = reset;
  assign mem_MPORT_462_data = 32'h0;
  assign mem_MPORT_462_addr = 9'h1ce;
  assign mem_MPORT_462_mask = 1'h1;
  assign mem_MPORT_462_en = reset;
  assign mem_MPORT_463_data = 32'h0;
  assign mem_MPORT_463_addr = 9'h1cf;
  assign mem_MPORT_463_mask = 1'h1;
  assign mem_MPORT_463_en = reset;
  assign mem_MPORT_464_data = 32'h0;
  assign mem_MPORT_464_addr = 9'h1d0;
  assign mem_MPORT_464_mask = 1'h1;
  assign mem_MPORT_464_en = reset;
  assign mem_MPORT_465_data = 32'h0;
  assign mem_MPORT_465_addr = 9'h1d1;
  assign mem_MPORT_465_mask = 1'h1;
  assign mem_MPORT_465_en = reset;
  assign mem_MPORT_466_data = 32'h0;
  assign mem_MPORT_466_addr = 9'h1d2;
  assign mem_MPORT_466_mask = 1'h1;
  assign mem_MPORT_466_en = reset;
  assign mem_MPORT_467_data = 32'h0;
  assign mem_MPORT_467_addr = 9'h1d3;
  assign mem_MPORT_467_mask = 1'h1;
  assign mem_MPORT_467_en = reset;
  assign mem_MPORT_468_data = 32'h0;
  assign mem_MPORT_468_addr = 9'h1d4;
  assign mem_MPORT_468_mask = 1'h1;
  assign mem_MPORT_468_en = reset;
  assign mem_MPORT_469_data = 32'h0;
  assign mem_MPORT_469_addr = 9'h1d5;
  assign mem_MPORT_469_mask = 1'h1;
  assign mem_MPORT_469_en = reset;
  assign mem_MPORT_470_data = 32'h0;
  assign mem_MPORT_470_addr = 9'h1d6;
  assign mem_MPORT_470_mask = 1'h1;
  assign mem_MPORT_470_en = reset;
  assign mem_MPORT_471_data = 32'h0;
  assign mem_MPORT_471_addr = 9'h1d7;
  assign mem_MPORT_471_mask = 1'h1;
  assign mem_MPORT_471_en = reset;
  assign mem_MPORT_472_data = 32'h0;
  assign mem_MPORT_472_addr = 9'h1d8;
  assign mem_MPORT_472_mask = 1'h1;
  assign mem_MPORT_472_en = reset;
  assign mem_MPORT_473_data = 32'h0;
  assign mem_MPORT_473_addr = 9'h1d9;
  assign mem_MPORT_473_mask = 1'h1;
  assign mem_MPORT_473_en = reset;
  assign mem_MPORT_474_data = 32'h0;
  assign mem_MPORT_474_addr = 9'h1da;
  assign mem_MPORT_474_mask = 1'h1;
  assign mem_MPORT_474_en = reset;
  assign mem_MPORT_475_data = 32'h0;
  assign mem_MPORT_475_addr = 9'h1db;
  assign mem_MPORT_475_mask = 1'h1;
  assign mem_MPORT_475_en = reset;
  assign mem_MPORT_476_data = 32'h0;
  assign mem_MPORT_476_addr = 9'h1dc;
  assign mem_MPORT_476_mask = 1'h1;
  assign mem_MPORT_476_en = reset;
  assign mem_MPORT_477_data = 32'h0;
  assign mem_MPORT_477_addr = 9'h1dd;
  assign mem_MPORT_477_mask = 1'h1;
  assign mem_MPORT_477_en = reset;
  assign mem_MPORT_478_data = 32'h0;
  assign mem_MPORT_478_addr = 9'h1de;
  assign mem_MPORT_478_mask = 1'h1;
  assign mem_MPORT_478_en = reset;
  assign mem_MPORT_479_data = 32'h0;
  assign mem_MPORT_479_addr = 9'h1df;
  assign mem_MPORT_479_mask = 1'h1;
  assign mem_MPORT_479_en = reset;
  assign mem_MPORT_480_data = 32'h0;
  assign mem_MPORT_480_addr = 9'h1e0;
  assign mem_MPORT_480_mask = 1'h1;
  assign mem_MPORT_480_en = reset;
  assign mem_MPORT_481_data = 32'h0;
  assign mem_MPORT_481_addr = 9'h1e1;
  assign mem_MPORT_481_mask = 1'h1;
  assign mem_MPORT_481_en = reset;
  assign mem_MPORT_482_data = 32'h0;
  assign mem_MPORT_482_addr = 9'h1e2;
  assign mem_MPORT_482_mask = 1'h1;
  assign mem_MPORT_482_en = reset;
  assign mem_MPORT_483_data = 32'h0;
  assign mem_MPORT_483_addr = 9'h1e3;
  assign mem_MPORT_483_mask = 1'h1;
  assign mem_MPORT_483_en = reset;
  assign mem_MPORT_484_data = 32'h0;
  assign mem_MPORT_484_addr = 9'h1e4;
  assign mem_MPORT_484_mask = 1'h1;
  assign mem_MPORT_484_en = reset;
  assign mem_MPORT_485_data = 32'h0;
  assign mem_MPORT_485_addr = 9'h1e5;
  assign mem_MPORT_485_mask = 1'h1;
  assign mem_MPORT_485_en = reset;
  assign mem_MPORT_486_data = 32'h0;
  assign mem_MPORT_486_addr = 9'h1e6;
  assign mem_MPORT_486_mask = 1'h1;
  assign mem_MPORT_486_en = reset;
  assign mem_MPORT_487_data = 32'h0;
  assign mem_MPORT_487_addr = 9'h1e7;
  assign mem_MPORT_487_mask = 1'h1;
  assign mem_MPORT_487_en = reset;
  assign mem_MPORT_488_data = 32'h0;
  assign mem_MPORT_488_addr = 9'h1e8;
  assign mem_MPORT_488_mask = 1'h1;
  assign mem_MPORT_488_en = reset;
  assign mem_MPORT_489_data = 32'h0;
  assign mem_MPORT_489_addr = 9'h1e9;
  assign mem_MPORT_489_mask = 1'h1;
  assign mem_MPORT_489_en = reset;
  assign mem_MPORT_490_data = 32'h0;
  assign mem_MPORT_490_addr = 9'h1ea;
  assign mem_MPORT_490_mask = 1'h1;
  assign mem_MPORT_490_en = reset;
  assign mem_MPORT_491_data = 32'h0;
  assign mem_MPORT_491_addr = 9'h1eb;
  assign mem_MPORT_491_mask = 1'h1;
  assign mem_MPORT_491_en = reset;
  assign mem_MPORT_492_data = 32'h0;
  assign mem_MPORT_492_addr = 9'h1ec;
  assign mem_MPORT_492_mask = 1'h1;
  assign mem_MPORT_492_en = reset;
  assign mem_MPORT_493_data = 32'h0;
  assign mem_MPORT_493_addr = 9'h1ed;
  assign mem_MPORT_493_mask = 1'h1;
  assign mem_MPORT_493_en = reset;
  assign mem_MPORT_494_data = 32'h0;
  assign mem_MPORT_494_addr = 9'h1ee;
  assign mem_MPORT_494_mask = 1'h1;
  assign mem_MPORT_494_en = reset;
  assign mem_MPORT_495_data = 32'h0;
  assign mem_MPORT_495_addr = 9'h1ef;
  assign mem_MPORT_495_mask = 1'h1;
  assign mem_MPORT_495_en = reset;
  assign mem_MPORT_496_data = 32'h0;
  assign mem_MPORT_496_addr = 9'h1f0;
  assign mem_MPORT_496_mask = 1'h1;
  assign mem_MPORT_496_en = reset;
  assign mem_MPORT_497_data = 32'h0;
  assign mem_MPORT_497_addr = 9'h1f1;
  assign mem_MPORT_497_mask = 1'h1;
  assign mem_MPORT_497_en = reset;
  assign mem_MPORT_498_data = 32'h0;
  assign mem_MPORT_498_addr = 9'h1f2;
  assign mem_MPORT_498_mask = 1'h1;
  assign mem_MPORT_498_en = reset;
  assign mem_MPORT_499_data = 32'h0;
  assign mem_MPORT_499_addr = 9'h1f3;
  assign mem_MPORT_499_mask = 1'h1;
  assign mem_MPORT_499_en = reset;
  assign mem_MPORT_500_data = 32'h0;
  assign mem_MPORT_500_addr = 9'h1f4;
  assign mem_MPORT_500_mask = 1'h1;
  assign mem_MPORT_500_en = reset;
  assign mem_MPORT_501_data = 32'h0;
  assign mem_MPORT_501_addr = 9'h1f5;
  assign mem_MPORT_501_mask = 1'h1;
  assign mem_MPORT_501_en = reset;
  assign mem_MPORT_502_data = 32'h0;
  assign mem_MPORT_502_addr = 9'h1f6;
  assign mem_MPORT_502_mask = 1'h1;
  assign mem_MPORT_502_en = reset;
  assign mem_MPORT_503_data = 32'h0;
  assign mem_MPORT_503_addr = 9'h1f7;
  assign mem_MPORT_503_mask = 1'h1;
  assign mem_MPORT_503_en = reset;
  assign mem_MPORT_504_data = 32'h0;
  assign mem_MPORT_504_addr = 9'h1f8;
  assign mem_MPORT_504_mask = 1'h1;
  assign mem_MPORT_504_en = reset;
  assign mem_MPORT_505_data = 32'h0;
  assign mem_MPORT_505_addr = 9'h1f9;
  assign mem_MPORT_505_mask = 1'h1;
  assign mem_MPORT_505_en = reset;
  assign mem_MPORT_506_data = 32'h0;
  assign mem_MPORT_506_addr = 9'h1fa;
  assign mem_MPORT_506_mask = 1'h1;
  assign mem_MPORT_506_en = reset;
  assign mem_MPORT_507_data = 32'h0;
  assign mem_MPORT_507_addr = 9'h1fb;
  assign mem_MPORT_507_mask = 1'h1;
  assign mem_MPORT_507_en = reset;
  assign mem_MPORT_508_data = 32'h0;
  assign mem_MPORT_508_addr = 9'h1fc;
  assign mem_MPORT_508_mask = 1'h1;
  assign mem_MPORT_508_en = reset;
  assign mem_MPORT_509_data = 32'h0;
  assign mem_MPORT_509_addr = 9'h1fd;
  assign mem_MPORT_509_mask = 1'h1;
  assign mem_MPORT_509_en = reset;
  assign mem_MPORT_510_data = 32'h0;
  assign mem_MPORT_510_addr = 9'h1fe;
  assign mem_MPORT_510_mask = 1'h1;
  assign mem_MPORT_510_en = reset;
  assign mem_MPORT_511_data = 32'h0;
  assign mem_MPORT_511_addr = 9'h1ff;
  assign mem_MPORT_511_mask = 1'h1;
  assign mem_MPORT_511_en = reset;
  assign mem_MPORT_512_data = io_w_data;
  assign mem_MPORT_512_addr = io_w_addr;
  assign mem_MPORT_512_mask = 1'h1;
  assign mem_MPORT_512_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_129_en & mem_MPORT_129_mask) begin
      mem[mem_MPORT_129_addr] <= mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_130_en & mem_MPORT_130_mask) begin
      mem[mem_MPORT_130_addr] <= mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_131_en & mem_MPORT_131_mask) begin
      mem[mem_MPORT_131_addr] <= mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_132_en & mem_MPORT_132_mask) begin
      mem[mem_MPORT_132_addr] <= mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_133_en & mem_MPORT_133_mask) begin
      mem[mem_MPORT_133_addr] <= mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_134_en & mem_MPORT_134_mask) begin
      mem[mem_MPORT_134_addr] <= mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_135_en & mem_MPORT_135_mask) begin
      mem[mem_MPORT_135_addr] <= mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_136_en & mem_MPORT_136_mask) begin
      mem[mem_MPORT_136_addr] <= mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_137_en & mem_MPORT_137_mask) begin
      mem[mem_MPORT_137_addr] <= mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_138_en & mem_MPORT_138_mask) begin
      mem[mem_MPORT_138_addr] <= mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_139_en & mem_MPORT_139_mask) begin
      mem[mem_MPORT_139_addr] <= mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_140_en & mem_MPORT_140_mask) begin
      mem[mem_MPORT_140_addr] <= mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_141_en & mem_MPORT_141_mask) begin
      mem[mem_MPORT_141_addr] <= mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_142_en & mem_MPORT_142_mask) begin
      mem[mem_MPORT_142_addr] <= mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_143_en & mem_MPORT_143_mask) begin
      mem[mem_MPORT_143_addr] <= mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_144_en & mem_MPORT_144_mask) begin
      mem[mem_MPORT_144_addr] <= mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_145_en & mem_MPORT_145_mask) begin
      mem[mem_MPORT_145_addr] <= mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_146_en & mem_MPORT_146_mask) begin
      mem[mem_MPORT_146_addr] <= mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_147_en & mem_MPORT_147_mask) begin
      mem[mem_MPORT_147_addr] <= mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_148_en & mem_MPORT_148_mask) begin
      mem[mem_MPORT_148_addr] <= mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_149_en & mem_MPORT_149_mask) begin
      mem[mem_MPORT_149_addr] <= mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_150_en & mem_MPORT_150_mask) begin
      mem[mem_MPORT_150_addr] <= mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_151_en & mem_MPORT_151_mask) begin
      mem[mem_MPORT_151_addr] <= mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_152_en & mem_MPORT_152_mask) begin
      mem[mem_MPORT_152_addr] <= mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_153_en & mem_MPORT_153_mask) begin
      mem[mem_MPORT_153_addr] <= mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_154_en & mem_MPORT_154_mask) begin
      mem[mem_MPORT_154_addr] <= mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_155_en & mem_MPORT_155_mask) begin
      mem[mem_MPORT_155_addr] <= mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_156_en & mem_MPORT_156_mask) begin
      mem[mem_MPORT_156_addr] <= mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_157_en & mem_MPORT_157_mask) begin
      mem[mem_MPORT_157_addr] <= mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_158_en & mem_MPORT_158_mask) begin
      mem[mem_MPORT_158_addr] <= mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_159_en & mem_MPORT_159_mask) begin
      mem[mem_MPORT_159_addr] <= mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_160_en & mem_MPORT_160_mask) begin
      mem[mem_MPORT_160_addr] <= mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_161_en & mem_MPORT_161_mask) begin
      mem[mem_MPORT_161_addr] <= mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_162_en & mem_MPORT_162_mask) begin
      mem[mem_MPORT_162_addr] <= mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_163_en & mem_MPORT_163_mask) begin
      mem[mem_MPORT_163_addr] <= mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_164_en & mem_MPORT_164_mask) begin
      mem[mem_MPORT_164_addr] <= mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_165_en & mem_MPORT_165_mask) begin
      mem[mem_MPORT_165_addr] <= mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_166_en & mem_MPORT_166_mask) begin
      mem[mem_MPORT_166_addr] <= mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_167_en & mem_MPORT_167_mask) begin
      mem[mem_MPORT_167_addr] <= mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_168_en & mem_MPORT_168_mask) begin
      mem[mem_MPORT_168_addr] <= mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_169_en & mem_MPORT_169_mask) begin
      mem[mem_MPORT_169_addr] <= mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_170_en & mem_MPORT_170_mask) begin
      mem[mem_MPORT_170_addr] <= mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_171_en & mem_MPORT_171_mask) begin
      mem[mem_MPORT_171_addr] <= mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_172_en & mem_MPORT_172_mask) begin
      mem[mem_MPORT_172_addr] <= mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_173_en & mem_MPORT_173_mask) begin
      mem[mem_MPORT_173_addr] <= mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_174_en & mem_MPORT_174_mask) begin
      mem[mem_MPORT_174_addr] <= mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_175_en & mem_MPORT_175_mask) begin
      mem[mem_MPORT_175_addr] <= mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_176_en & mem_MPORT_176_mask) begin
      mem[mem_MPORT_176_addr] <= mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_177_en & mem_MPORT_177_mask) begin
      mem[mem_MPORT_177_addr] <= mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_178_en & mem_MPORT_178_mask) begin
      mem[mem_MPORT_178_addr] <= mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_179_en & mem_MPORT_179_mask) begin
      mem[mem_MPORT_179_addr] <= mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_180_en & mem_MPORT_180_mask) begin
      mem[mem_MPORT_180_addr] <= mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_181_en & mem_MPORT_181_mask) begin
      mem[mem_MPORT_181_addr] <= mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_182_en & mem_MPORT_182_mask) begin
      mem[mem_MPORT_182_addr] <= mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_183_en & mem_MPORT_183_mask) begin
      mem[mem_MPORT_183_addr] <= mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_184_en & mem_MPORT_184_mask) begin
      mem[mem_MPORT_184_addr] <= mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_185_en & mem_MPORT_185_mask) begin
      mem[mem_MPORT_185_addr] <= mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_186_en & mem_MPORT_186_mask) begin
      mem[mem_MPORT_186_addr] <= mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_187_en & mem_MPORT_187_mask) begin
      mem[mem_MPORT_187_addr] <= mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_188_en & mem_MPORT_188_mask) begin
      mem[mem_MPORT_188_addr] <= mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_189_en & mem_MPORT_189_mask) begin
      mem[mem_MPORT_189_addr] <= mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_190_en & mem_MPORT_190_mask) begin
      mem[mem_MPORT_190_addr] <= mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_191_en & mem_MPORT_191_mask) begin
      mem[mem_MPORT_191_addr] <= mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_192_en & mem_MPORT_192_mask) begin
      mem[mem_MPORT_192_addr] <= mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_193_en & mem_MPORT_193_mask) begin
      mem[mem_MPORT_193_addr] <= mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_194_en & mem_MPORT_194_mask) begin
      mem[mem_MPORT_194_addr] <= mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_195_en & mem_MPORT_195_mask) begin
      mem[mem_MPORT_195_addr] <= mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_196_en & mem_MPORT_196_mask) begin
      mem[mem_MPORT_196_addr] <= mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_197_en & mem_MPORT_197_mask) begin
      mem[mem_MPORT_197_addr] <= mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_198_en & mem_MPORT_198_mask) begin
      mem[mem_MPORT_198_addr] <= mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_199_en & mem_MPORT_199_mask) begin
      mem[mem_MPORT_199_addr] <= mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_200_en & mem_MPORT_200_mask) begin
      mem[mem_MPORT_200_addr] <= mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_201_en & mem_MPORT_201_mask) begin
      mem[mem_MPORT_201_addr] <= mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_202_en & mem_MPORT_202_mask) begin
      mem[mem_MPORT_202_addr] <= mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_203_en & mem_MPORT_203_mask) begin
      mem[mem_MPORT_203_addr] <= mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_204_en & mem_MPORT_204_mask) begin
      mem[mem_MPORT_204_addr] <= mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_205_en & mem_MPORT_205_mask) begin
      mem[mem_MPORT_205_addr] <= mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_206_en & mem_MPORT_206_mask) begin
      mem[mem_MPORT_206_addr] <= mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_207_en & mem_MPORT_207_mask) begin
      mem[mem_MPORT_207_addr] <= mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_208_en & mem_MPORT_208_mask) begin
      mem[mem_MPORT_208_addr] <= mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_209_en & mem_MPORT_209_mask) begin
      mem[mem_MPORT_209_addr] <= mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_210_en & mem_MPORT_210_mask) begin
      mem[mem_MPORT_210_addr] <= mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_211_en & mem_MPORT_211_mask) begin
      mem[mem_MPORT_211_addr] <= mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_212_en & mem_MPORT_212_mask) begin
      mem[mem_MPORT_212_addr] <= mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_213_en & mem_MPORT_213_mask) begin
      mem[mem_MPORT_213_addr] <= mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_214_en & mem_MPORT_214_mask) begin
      mem[mem_MPORT_214_addr] <= mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_215_en & mem_MPORT_215_mask) begin
      mem[mem_MPORT_215_addr] <= mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_216_en & mem_MPORT_216_mask) begin
      mem[mem_MPORT_216_addr] <= mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_217_en & mem_MPORT_217_mask) begin
      mem[mem_MPORT_217_addr] <= mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_218_en & mem_MPORT_218_mask) begin
      mem[mem_MPORT_218_addr] <= mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_219_en & mem_MPORT_219_mask) begin
      mem[mem_MPORT_219_addr] <= mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_220_en & mem_MPORT_220_mask) begin
      mem[mem_MPORT_220_addr] <= mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_221_en & mem_MPORT_221_mask) begin
      mem[mem_MPORT_221_addr] <= mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_222_en & mem_MPORT_222_mask) begin
      mem[mem_MPORT_222_addr] <= mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_223_en & mem_MPORT_223_mask) begin
      mem[mem_MPORT_223_addr] <= mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_224_en & mem_MPORT_224_mask) begin
      mem[mem_MPORT_224_addr] <= mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_225_en & mem_MPORT_225_mask) begin
      mem[mem_MPORT_225_addr] <= mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_226_en & mem_MPORT_226_mask) begin
      mem[mem_MPORT_226_addr] <= mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_227_en & mem_MPORT_227_mask) begin
      mem[mem_MPORT_227_addr] <= mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_228_en & mem_MPORT_228_mask) begin
      mem[mem_MPORT_228_addr] <= mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_229_en & mem_MPORT_229_mask) begin
      mem[mem_MPORT_229_addr] <= mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_230_en & mem_MPORT_230_mask) begin
      mem[mem_MPORT_230_addr] <= mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_231_en & mem_MPORT_231_mask) begin
      mem[mem_MPORT_231_addr] <= mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_232_en & mem_MPORT_232_mask) begin
      mem[mem_MPORT_232_addr] <= mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_233_en & mem_MPORT_233_mask) begin
      mem[mem_MPORT_233_addr] <= mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_234_en & mem_MPORT_234_mask) begin
      mem[mem_MPORT_234_addr] <= mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_235_en & mem_MPORT_235_mask) begin
      mem[mem_MPORT_235_addr] <= mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_236_en & mem_MPORT_236_mask) begin
      mem[mem_MPORT_236_addr] <= mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_237_en & mem_MPORT_237_mask) begin
      mem[mem_MPORT_237_addr] <= mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_238_en & mem_MPORT_238_mask) begin
      mem[mem_MPORT_238_addr] <= mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_239_en & mem_MPORT_239_mask) begin
      mem[mem_MPORT_239_addr] <= mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_240_en & mem_MPORT_240_mask) begin
      mem[mem_MPORT_240_addr] <= mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_241_en & mem_MPORT_241_mask) begin
      mem[mem_MPORT_241_addr] <= mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_242_en & mem_MPORT_242_mask) begin
      mem[mem_MPORT_242_addr] <= mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_243_en & mem_MPORT_243_mask) begin
      mem[mem_MPORT_243_addr] <= mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_244_en & mem_MPORT_244_mask) begin
      mem[mem_MPORT_244_addr] <= mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_245_en & mem_MPORT_245_mask) begin
      mem[mem_MPORT_245_addr] <= mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_246_en & mem_MPORT_246_mask) begin
      mem[mem_MPORT_246_addr] <= mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_247_en & mem_MPORT_247_mask) begin
      mem[mem_MPORT_247_addr] <= mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_248_en & mem_MPORT_248_mask) begin
      mem[mem_MPORT_248_addr] <= mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_249_en & mem_MPORT_249_mask) begin
      mem[mem_MPORT_249_addr] <= mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_250_en & mem_MPORT_250_mask) begin
      mem[mem_MPORT_250_addr] <= mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_251_en & mem_MPORT_251_mask) begin
      mem[mem_MPORT_251_addr] <= mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_252_en & mem_MPORT_252_mask) begin
      mem[mem_MPORT_252_addr] <= mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_253_en & mem_MPORT_253_mask) begin
      mem[mem_MPORT_253_addr] <= mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_254_en & mem_MPORT_254_mask) begin
      mem[mem_MPORT_254_addr] <= mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_255_en & mem_MPORT_255_mask) begin
      mem[mem_MPORT_255_addr] <= mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_256_en & mem_MPORT_256_mask) begin
      mem[mem_MPORT_256_addr] <= mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_257_en & mem_MPORT_257_mask) begin
      mem[mem_MPORT_257_addr] <= mem_MPORT_257_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_258_en & mem_MPORT_258_mask) begin
      mem[mem_MPORT_258_addr] <= mem_MPORT_258_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_259_en & mem_MPORT_259_mask) begin
      mem[mem_MPORT_259_addr] <= mem_MPORT_259_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_260_en & mem_MPORT_260_mask) begin
      mem[mem_MPORT_260_addr] <= mem_MPORT_260_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_261_en & mem_MPORT_261_mask) begin
      mem[mem_MPORT_261_addr] <= mem_MPORT_261_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_262_en & mem_MPORT_262_mask) begin
      mem[mem_MPORT_262_addr] <= mem_MPORT_262_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_263_en & mem_MPORT_263_mask) begin
      mem[mem_MPORT_263_addr] <= mem_MPORT_263_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_264_en & mem_MPORT_264_mask) begin
      mem[mem_MPORT_264_addr] <= mem_MPORT_264_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_265_en & mem_MPORT_265_mask) begin
      mem[mem_MPORT_265_addr] <= mem_MPORT_265_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_266_en & mem_MPORT_266_mask) begin
      mem[mem_MPORT_266_addr] <= mem_MPORT_266_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_267_en & mem_MPORT_267_mask) begin
      mem[mem_MPORT_267_addr] <= mem_MPORT_267_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_268_en & mem_MPORT_268_mask) begin
      mem[mem_MPORT_268_addr] <= mem_MPORT_268_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_269_en & mem_MPORT_269_mask) begin
      mem[mem_MPORT_269_addr] <= mem_MPORT_269_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_270_en & mem_MPORT_270_mask) begin
      mem[mem_MPORT_270_addr] <= mem_MPORT_270_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_271_en & mem_MPORT_271_mask) begin
      mem[mem_MPORT_271_addr] <= mem_MPORT_271_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_272_en & mem_MPORT_272_mask) begin
      mem[mem_MPORT_272_addr] <= mem_MPORT_272_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_273_en & mem_MPORT_273_mask) begin
      mem[mem_MPORT_273_addr] <= mem_MPORT_273_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_274_en & mem_MPORT_274_mask) begin
      mem[mem_MPORT_274_addr] <= mem_MPORT_274_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_275_en & mem_MPORT_275_mask) begin
      mem[mem_MPORT_275_addr] <= mem_MPORT_275_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_276_en & mem_MPORT_276_mask) begin
      mem[mem_MPORT_276_addr] <= mem_MPORT_276_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_277_en & mem_MPORT_277_mask) begin
      mem[mem_MPORT_277_addr] <= mem_MPORT_277_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_278_en & mem_MPORT_278_mask) begin
      mem[mem_MPORT_278_addr] <= mem_MPORT_278_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_279_en & mem_MPORT_279_mask) begin
      mem[mem_MPORT_279_addr] <= mem_MPORT_279_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_280_en & mem_MPORT_280_mask) begin
      mem[mem_MPORT_280_addr] <= mem_MPORT_280_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_281_en & mem_MPORT_281_mask) begin
      mem[mem_MPORT_281_addr] <= mem_MPORT_281_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_282_en & mem_MPORT_282_mask) begin
      mem[mem_MPORT_282_addr] <= mem_MPORT_282_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_283_en & mem_MPORT_283_mask) begin
      mem[mem_MPORT_283_addr] <= mem_MPORT_283_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_284_en & mem_MPORT_284_mask) begin
      mem[mem_MPORT_284_addr] <= mem_MPORT_284_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_285_en & mem_MPORT_285_mask) begin
      mem[mem_MPORT_285_addr] <= mem_MPORT_285_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_286_en & mem_MPORT_286_mask) begin
      mem[mem_MPORT_286_addr] <= mem_MPORT_286_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_287_en & mem_MPORT_287_mask) begin
      mem[mem_MPORT_287_addr] <= mem_MPORT_287_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_288_en & mem_MPORT_288_mask) begin
      mem[mem_MPORT_288_addr] <= mem_MPORT_288_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_289_en & mem_MPORT_289_mask) begin
      mem[mem_MPORT_289_addr] <= mem_MPORT_289_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_290_en & mem_MPORT_290_mask) begin
      mem[mem_MPORT_290_addr] <= mem_MPORT_290_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_291_en & mem_MPORT_291_mask) begin
      mem[mem_MPORT_291_addr] <= mem_MPORT_291_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_292_en & mem_MPORT_292_mask) begin
      mem[mem_MPORT_292_addr] <= mem_MPORT_292_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_293_en & mem_MPORT_293_mask) begin
      mem[mem_MPORT_293_addr] <= mem_MPORT_293_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_294_en & mem_MPORT_294_mask) begin
      mem[mem_MPORT_294_addr] <= mem_MPORT_294_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_295_en & mem_MPORT_295_mask) begin
      mem[mem_MPORT_295_addr] <= mem_MPORT_295_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_296_en & mem_MPORT_296_mask) begin
      mem[mem_MPORT_296_addr] <= mem_MPORT_296_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_297_en & mem_MPORT_297_mask) begin
      mem[mem_MPORT_297_addr] <= mem_MPORT_297_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_298_en & mem_MPORT_298_mask) begin
      mem[mem_MPORT_298_addr] <= mem_MPORT_298_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_299_en & mem_MPORT_299_mask) begin
      mem[mem_MPORT_299_addr] <= mem_MPORT_299_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_300_en & mem_MPORT_300_mask) begin
      mem[mem_MPORT_300_addr] <= mem_MPORT_300_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_301_en & mem_MPORT_301_mask) begin
      mem[mem_MPORT_301_addr] <= mem_MPORT_301_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_302_en & mem_MPORT_302_mask) begin
      mem[mem_MPORT_302_addr] <= mem_MPORT_302_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_303_en & mem_MPORT_303_mask) begin
      mem[mem_MPORT_303_addr] <= mem_MPORT_303_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_304_en & mem_MPORT_304_mask) begin
      mem[mem_MPORT_304_addr] <= mem_MPORT_304_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_305_en & mem_MPORT_305_mask) begin
      mem[mem_MPORT_305_addr] <= mem_MPORT_305_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_306_en & mem_MPORT_306_mask) begin
      mem[mem_MPORT_306_addr] <= mem_MPORT_306_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_307_en & mem_MPORT_307_mask) begin
      mem[mem_MPORT_307_addr] <= mem_MPORT_307_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_308_en & mem_MPORT_308_mask) begin
      mem[mem_MPORT_308_addr] <= mem_MPORT_308_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_309_en & mem_MPORT_309_mask) begin
      mem[mem_MPORT_309_addr] <= mem_MPORT_309_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_310_en & mem_MPORT_310_mask) begin
      mem[mem_MPORT_310_addr] <= mem_MPORT_310_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_311_en & mem_MPORT_311_mask) begin
      mem[mem_MPORT_311_addr] <= mem_MPORT_311_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_312_en & mem_MPORT_312_mask) begin
      mem[mem_MPORT_312_addr] <= mem_MPORT_312_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_313_en & mem_MPORT_313_mask) begin
      mem[mem_MPORT_313_addr] <= mem_MPORT_313_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_314_en & mem_MPORT_314_mask) begin
      mem[mem_MPORT_314_addr] <= mem_MPORT_314_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_315_en & mem_MPORT_315_mask) begin
      mem[mem_MPORT_315_addr] <= mem_MPORT_315_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_316_en & mem_MPORT_316_mask) begin
      mem[mem_MPORT_316_addr] <= mem_MPORT_316_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_317_en & mem_MPORT_317_mask) begin
      mem[mem_MPORT_317_addr] <= mem_MPORT_317_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_318_en & mem_MPORT_318_mask) begin
      mem[mem_MPORT_318_addr] <= mem_MPORT_318_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_319_en & mem_MPORT_319_mask) begin
      mem[mem_MPORT_319_addr] <= mem_MPORT_319_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_320_en & mem_MPORT_320_mask) begin
      mem[mem_MPORT_320_addr] <= mem_MPORT_320_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_321_en & mem_MPORT_321_mask) begin
      mem[mem_MPORT_321_addr] <= mem_MPORT_321_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_322_en & mem_MPORT_322_mask) begin
      mem[mem_MPORT_322_addr] <= mem_MPORT_322_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_323_en & mem_MPORT_323_mask) begin
      mem[mem_MPORT_323_addr] <= mem_MPORT_323_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_324_en & mem_MPORT_324_mask) begin
      mem[mem_MPORT_324_addr] <= mem_MPORT_324_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_325_en & mem_MPORT_325_mask) begin
      mem[mem_MPORT_325_addr] <= mem_MPORT_325_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_326_en & mem_MPORT_326_mask) begin
      mem[mem_MPORT_326_addr] <= mem_MPORT_326_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_327_en & mem_MPORT_327_mask) begin
      mem[mem_MPORT_327_addr] <= mem_MPORT_327_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_328_en & mem_MPORT_328_mask) begin
      mem[mem_MPORT_328_addr] <= mem_MPORT_328_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_329_en & mem_MPORT_329_mask) begin
      mem[mem_MPORT_329_addr] <= mem_MPORT_329_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_330_en & mem_MPORT_330_mask) begin
      mem[mem_MPORT_330_addr] <= mem_MPORT_330_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_331_en & mem_MPORT_331_mask) begin
      mem[mem_MPORT_331_addr] <= mem_MPORT_331_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_332_en & mem_MPORT_332_mask) begin
      mem[mem_MPORT_332_addr] <= mem_MPORT_332_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_333_en & mem_MPORT_333_mask) begin
      mem[mem_MPORT_333_addr] <= mem_MPORT_333_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_334_en & mem_MPORT_334_mask) begin
      mem[mem_MPORT_334_addr] <= mem_MPORT_334_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_335_en & mem_MPORT_335_mask) begin
      mem[mem_MPORT_335_addr] <= mem_MPORT_335_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_336_en & mem_MPORT_336_mask) begin
      mem[mem_MPORT_336_addr] <= mem_MPORT_336_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_337_en & mem_MPORT_337_mask) begin
      mem[mem_MPORT_337_addr] <= mem_MPORT_337_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_338_en & mem_MPORT_338_mask) begin
      mem[mem_MPORT_338_addr] <= mem_MPORT_338_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_339_en & mem_MPORT_339_mask) begin
      mem[mem_MPORT_339_addr] <= mem_MPORT_339_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_340_en & mem_MPORT_340_mask) begin
      mem[mem_MPORT_340_addr] <= mem_MPORT_340_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_341_en & mem_MPORT_341_mask) begin
      mem[mem_MPORT_341_addr] <= mem_MPORT_341_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_342_en & mem_MPORT_342_mask) begin
      mem[mem_MPORT_342_addr] <= mem_MPORT_342_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_343_en & mem_MPORT_343_mask) begin
      mem[mem_MPORT_343_addr] <= mem_MPORT_343_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_344_en & mem_MPORT_344_mask) begin
      mem[mem_MPORT_344_addr] <= mem_MPORT_344_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_345_en & mem_MPORT_345_mask) begin
      mem[mem_MPORT_345_addr] <= mem_MPORT_345_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_346_en & mem_MPORT_346_mask) begin
      mem[mem_MPORT_346_addr] <= mem_MPORT_346_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_347_en & mem_MPORT_347_mask) begin
      mem[mem_MPORT_347_addr] <= mem_MPORT_347_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_348_en & mem_MPORT_348_mask) begin
      mem[mem_MPORT_348_addr] <= mem_MPORT_348_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_349_en & mem_MPORT_349_mask) begin
      mem[mem_MPORT_349_addr] <= mem_MPORT_349_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_350_en & mem_MPORT_350_mask) begin
      mem[mem_MPORT_350_addr] <= mem_MPORT_350_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_351_en & mem_MPORT_351_mask) begin
      mem[mem_MPORT_351_addr] <= mem_MPORT_351_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_352_en & mem_MPORT_352_mask) begin
      mem[mem_MPORT_352_addr] <= mem_MPORT_352_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_353_en & mem_MPORT_353_mask) begin
      mem[mem_MPORT_353_addr] <= mem_MPORT_353_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_354_en & mem_MPORT_354_mask) begin
      mem[mem_MPORT_354_addr] <= mem_MPORT_354_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_355_en & mem_MPORT_355_mask) begin
      mem[mem_MPORT_355_addr] <= mem_MPORT_355_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_356_en & mem_MPORT_356_mask) begin
      mem[mem_MPORT_356_addr] <= mem_MPORT_356_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_357_en & mem_MPORT_357_mask) begin
      mem[mem_MPORT_357_addr] <= mem_MPORT_357_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_358_en & mem_MPORT_358_mask) begin
      mem[mem_MPORT_358_addr] <= mem_MPORT_358_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_359_en & mem_MPORT_359_mask) begin
      mem[mem_MPORT_359_addr] <= mem_MPORT_359_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_360_en & mem_MPORT_360_mask) begin
      mem[mem_MPORT_360_addr] <= mem_MPORT_360_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_361_en & mem_MPORT_361_mask) begin
      mem[mem_MPORT_361_addr] <= mem_MPORT_361_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_362_en & mem_MPORT_362_mask) begin
      mem[mem_MPORT_362_addr] <= mem_MPORT_362_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_363_en & mem_MPORT_363_mask) begin
      mem[mem_MPORT_363_addr] <= mem_MPORT_363_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_364_en & mem_MPORT_364_mask) begin
      mem[mem_MPORT_364_addr] <= mem_MPORT_364_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_365_en & mem_MPORT_365_mask) begin
      mem[mem_MPORT_365_addr] <= mem_MPORT_365_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_366_en & mem_MPORT_366_mask) begin
      mem[mem_MPORT_366_addr] <= mem_MPORT_366_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_367_en & mem_MPORT_367_mask) begin
      mem[mem_MPORT_367_addr] <= mem_MPORT_367_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_368_en & mem_MPORT_368_mask) begin
      mem[mem_MPORT_368_addr] <= mem_MPORT_368_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_369_en & mem_MPORT_369_mask) begin
      mem[mem_MPORT_369_addr] <= mem_MPORT_369_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_370_en & mem_MPORT_370_mask) begin
      mem[mem_MPORT_370_addr] <= mem_MPORT_370_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_371_en & mem_MPORT_371_mask) begin
      mem[mem_MPORT_371_addr] <= mem_MPORT_371_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_372_en & mem_MPORT_372_mask) begin
      mem[mem_MPORT_372_addr] <= mem_MPORT_372_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_373_en & mem_MPORT_373_mask) begin
      mem[mem_MPORT_373_addr] <= mem_MPORT_373_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_374_en & mem_MPORT_374_mask) begin
      mem[mem_MPORT_374_addr] <= mem_MPORT_374_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_375_en & mem_MPORT_375_mask) begin
      mem[mem_MPORT_375_addr] <= mem_MPORT_375_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_376_en & mem_MPORT_376_mask) begin
      mem[mem_MPORT_376_addr] <= mem_MPORT_376_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_377_en & mem_MPORT_377_mask) begin
      mem[mem_MPORT_377_addr] <= mem_MPORT_377_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_378_en & mem_MPORT_378_mask) begin
      mem[mem_MPORT_378_addr] <= mem_MPORT_378_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_379_en & mem_MPORT_379_mask) begin
      mem[mem_MPORT_379_addr] <= mem_MPORT_379_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_380_en & mem_MPORT_380_mask) begin
      mem[mem_MPORT_380_addr] <= mem_MPORT_380_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_381_en & mem_MPORT_381_mask) begin
      mem[mem_MPORT_381_addr] <= mem_MPORT_381_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_382_en & mem_MPORT_382_mask) begin
      mem[mem_MPORT_382_addr] <= mem_MPORT_382_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_383_en & mem_MPORT_383_mask) begin
      mem[mem_MPORT_383_addr] <= mem_MPORT_383_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_384_en & mem_MPORT_384_mask) begin
      mem[mem_MPORT_384_addr] <= mem_MPORT_384_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_385_en & mem_MPORT_385_mask) begin
      mem[mem_MPORT_385_addr] <= mem_MPORT_385_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_386_en & mem_MPORT_386_mask) begin
      mem[mem_MPORT_386_addr] <= mem_MPORT_386_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_387_en & mem_MPORT_387_mask) begin
      mem[mem_MPORT_387_addr] <= mem_MPORT_387_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_388_en & mem_MPORT_388_mask) begin
      mem[mem_MPORT_388_addr] <= mem_MPORT_388_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_389_en & mem_MPORT_389_mask) begin
      mem[mem_MPORT_389_addr] <= mem_MPORT_389_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_390_en & mem_MPORT_390_mask) begin
      mem[mem_MPORT_390_addr] <= mem_MPORT_390_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_391_en & mem_MPORT_391_mask) begin
      mem[mem_MPORT_391_addr] <= mem_MPORT_391_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_392_en & mem_MPORT_392_mask) begin
      mem[mem_MPORT_392_addr] <= mem_MPORT_392_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_393_en & mem_MPORT_393_mask) begin
      mem[mem_MPORT_393_addr] <= mem_MPORT_393_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_394_en & mem_MPORT_394_mask) begin
      mem[mem_MPORT_394_addr] <= mem_MPORT_394_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_395_en & mem_MPORT_395_mask) begin
      mem[mem_MPORT_395_addr] <= mem_MPORT_395_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_396_en & mem_MPORT_396_mask) begin
      mem[mem_MPORT_396_addr] <= mem_MPORT_396_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_397_en & mem_MPORT_397_mask) begin
      mem[mem_MPORT_397_addr] <= mem_MPORT_397_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_398_en & mem_MPORT_398_mask) begin
      mem[mem_MPORT_398_addr] <= mem_MPORT_398_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_399_en & mem_MPORT_399_mask) begin
      mem[mem_MPORT_399_addr] <= mem_MPORT_399_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_400_en & mem_MPORT_400_mask) begin
      mem[mem_MPORT_400_addr] <= mem_MPORT_400_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_401_en & mem_MPORT_401_mask) begin
      mem[mem_MPORT_401_addr] <= mem_MPORT_401_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_402_en & mem_MPORT_402_mask) begin
      mem[mem_MPORT_402_addr] <= mem_MPORT_402_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_403_en & mem_MPORT_403_mask) begin
      mem[mem_MPORT_403_addr] <= mem_MPORT_403_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_404_en & mem_MPORT_404_mask) begin
      mem[mem_MPORT_404_addr] <= mem_MPORT_404_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_405_en & mem_MPORT_405_mask) begin
      mem[mem_MPORT_405_addr] <= mem_MPORT_405_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_406_en & mem_MPORT_406_mask) begin
      mem[mem_MPORT_406_addr] <= mem_MPORT_406_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_407_en & mem_MPORT_407_mask) begin
      mem[mem_MPORT_407_addr] <= mem_MPORT_407_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_408_en & mem_MPORT_408_mask) begin
      mem[mem_MPORT_408_addr] <= mem_MPORT_408_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_409_en & mem_MPORT_409_mask) begin
      mem[mem_MPORT_409_addr] <= mem_MPORT_409_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_410_en & mem_MPORT_410_mask) begin
      mem[mem_MPORT_410_addr] <= mem_MPORT_410_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_411_en & mem_MPORT_411_mask) begin
      mem[mem_MPORT_411_addr] <= mem_MPORT_411_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_412_en & mem_MPORT_412_mask) begin
      mem[mem_MPORT_412_addr] <= mem_MPORT_412_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_413_en & mem_MPORT_413_mask) begin
      mem[mem_MPORT_413_addr] <= mem_MPORT_413_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_414_en & mem_MPORT_414_mask) begin
      mem[mem_MPORT_414_addr] <= mem_MPORT_414_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_415_en & mem_MPORT_415_mask) begin
      mem[mem_MPORT_415_addr] <= mem_MPORT_415_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_416_en & mem_MPORT_416_mask) begin
      mem[mem_MPORT_416_addr] <= mem_MPORT_416_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_417_en & mem_MPORT_417_mask) begin
      mem[mem_MPORT_417_addr] <= mem_MPORT_417_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_418_en & mem_MPORT_418_mask) begin
      mem[mem_MPORT_418_addr] <= mem_MPORT_418_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_419_en & mem_MPORT_419_mask) begin
      mem[mem_MPORT_419_addr] <= mem_MPORT_419_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_420_en & mem_MPORT_420_mask) begin
      mem[mem_MPORT_420_addr] <= mem_MPORT_420_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_421_en & mem_MPORT_421_mask) begin
      mem[mem_MPORT_421_addr] <= mem_MPORT_421_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_422_en & mem_MPORT_422_mask) begin
      mem[mem_MPORT_422_addr] <= mem_MPORT_422_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_423_en & mem_MPORT_423_mask) begin
      mem[mem_MPORT_423_addr] <= mem_MPORT_423_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_424_en & mem_MPORT_424_mask) begin
      mem[mem_MPORT_424_addr] <= mem_MPORT_424_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_425_en & mem_MPORT_425_mask) begin
      mem[mem_MPORT_425_addr] <= mem_MPORT_425_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_426_en & mem_MPORT_426_mask) begin
      mem[mem_MPORT_426_addr] <= mem_MPORT_426_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_427_en & mem_MPORT_427_mask) begin
      mem[mem_MPORT_427_addr] <= mem_MPORT_427_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_428_en & mem_MPORT_428_mask) begin
      mem[mem_MPORT_428_addr] <= mem_MPORT_428_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_429_en & mem_MPORT_429_mask) begin
      mem[mem_MPORT_429_addr] <= mem_MPORT_429_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_430_en & mem_MPORT_430_mask) begin
      mem[mem_MPORT_430_addr] <= mem_MPORT_430_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_431_en & mem_MPORT_431_mask) begin
      mem[mem_MPORT_431_addr] <= mem_MPORT_431_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_432_en & mem_MPORT_432_mask) begin
      mem[mem_MPORT_432_addr] <= mem_MPORT_432_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_433_en & mem_MPORT_433_mask) begin
      mem[mem_MPORT_433_addr] <= mem_MPORT_433_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_434_en & mem_MPORT_434_mask) begin
      mem[mem_MPORT_434_addr] <= mem_MPORT_434_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_435_en & mem_MPORT_435_mask) begin
      mem[mem_MPORT_435_addr] <= mem_MPORT_435_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_436_en & mem_MPORT_436_mask) begin
      mem[mem_MPORT_436_addr] <= mem_MPORT_436_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_437_en & mem_MPORT_437_mask) begin
      mem[mem_MPORT_437_addr] <= mem_MPORT_437_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_438_en & mem_MPORT_438_mask) begin
      mem[mem_MPORT_438_addr] <= mem_MPORT_438_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_439_en & mem_MPORT_439_mask) begin
      mem[mem_MPORT_439_addr] <= mem_MPORT_439_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_440_en & mem_MPORT_440_mask) begin
      mem[mem_MPORT_440_addr] <= mem_MPORT_440_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_441_en & mem_MPORT_441_mask) begin
      mem[mem_MPORT_441_addr] <= mem_MPORT_441_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_442_en & mem_MPORT_442_mask) begin
      mem[mem_MPORT_442_addr] <= mem_MPORT_442_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_443_en & mem_MPORT_443_mask) begin
      mem[mem_MPORT_443_addr] <= mem_MPORT_443_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_444_en & mem_MPORT_444_mask) begin
      mem[mem_MPORT_444_addr] <= mem_MPORT_444_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_445_en & mem_MPORT_445_mask) begin
      mem[mem_MPORT_445_addr] <= mem_MPORT_445_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_446_en & mem_MPORT_446_mask) begin
      mem[mem_MPORT_446_addr] <= mem_MPORT_446_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_447_en & mem_MPORT_447_mask) begin
      mem[mem_MPORT_447_addr] <= mem_MPORT_447_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_448_en & mem_MPORT_448_mask) begin
      mem[mem_MPORT_448_addr] <= mem_MPORT_448_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_449_en & mem_MPORT_449_mask) begin
      mem[mem_MPORT_449_addr] <= mem_MPORT_449_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_450_en & mem_MPORT_450_mask) begin
      mem[mem_MPORT_450_addr] <= mem_MPORT_450_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_451_en & mem_MPORT_451_mask) begin
      mem[mem_MPORT_451_addr] <= mem_MPORT_451_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_452_en & mem_MPORT_452_mask) begin
      mem[mem_MPORT_452_addr] <= mem_MPORT_452_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_453_en & mem_MPORT_453_mask) begin
      mem[mem_MPORT_453_addr] <= mem_MPORT_453_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_454_en & mem_MPORT_454_mask) begin
      mem[mem_MPORT_454_addr] <= mem_MPORT_454_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_455_en & mem_MPORT_455_mask) begin
      mem[mem_MPORT_455_addr] <= mem_MPORT_455_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_456_en & mem_MPORT_456_mask) begin
      mem[mem_MPORT_456_addr] <= mem_MPORT_456_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_457_en & mem_MPORT_457_mask) begin
      mem[mem_MPORT_457_addr] <= mem_MPORT_457_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_458_en & mem_MPORT_458_mask) begin
      mem[mem_MPORT_458_addr] <= mem_MPORT_458_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_459_en & mem_MPORT_459_mask) begin
      mem[mem_MPORT_459_addr] <= mem_MPORT_459_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_460_en & mem_MPORT_460_mask) begin
      mem[mem_MPORT_460_addr] <= mem_MPORT_460_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_461_en & mem_MPORT_461_mask) begin
      mem[mem_MPORT_461_addr] <= mem_MPORT_461_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_462_en & mem_MPORT_462_mask) begin
      mem[mem_MPORT_462_addr] <= mem_MPORT_462_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_463_en & mem_MPORT_463_mask) begin
      mem[mem_MPORT_463_addr] <= mem_MPORT_463_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_464_en & mem_MPORT_464_mask) begin
      mem[mem_MPORT_464_addr] <= mem_MPORT_464_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_465_en & mem_MPORT_465_mask) begin
      mem[mem_MPORT_465_addr] <= mem_MPORT_465_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_466_en & mem_MPORT_466_mask) begin
      mem[mem_MPORT_466_addr] <= mem_MPORT_466_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_467_en & mem_MPORT_467_mask) begin
      mem[mem_MPORT_467_addr] <= mem_MPORT_467_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_468_en & mem_MPORT_468_mask) begin
      mem[mem_MPORT_468_addr] <= mem_MPORT_468_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_469_en & mem_MPORT_469_mask) begin
      mem[mem_MPORT_469_addr] <= mem_MPORT_469_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_470_en & mem_MPORT_470_mask) begin
      mem[mem_MPORT_470_addr] <= mem_MPORT_470_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_471_en & mem_MPORT_471_mask) begin
      mem[mem_MPORT_471_addr] <= mem_MPORT_471_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_472_en & mem_MPORT_472_mask) begin
      mem[mem_MPORT_472_addr] <= mem_MPORT_472_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_473_en & mem_MPORT_473_mask) begin
      mem[mem_MPORT_473_addr] <= mem_MPORT_473_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_474_en & mem_MPORT_474_mask) begin
      mem[mem_MPORT_474_addr] <= mem_MPORT_474_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_475_en & mem_MPORT_475_mask) begin
      mem[mem_MPORT_475_addr] <= mem_MPORT_475_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_476_en & mem_MPORT_476_mask) begin
      mem[mem_MPORT_476_addr] <= mem_MPORT_476_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_477_en & mem_MPORT_477_mask) begin
      mem[mem_MPORT_477_addr] <= mem_MPORT_477_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_478_en & mem_MPORT_478_mask) begin
      mem[mem_MPORT_478_addr] <= mem_MPORT_478_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_479_en & mem_MPORT_479_mask) begin
      mem[mem_MPORT_479_addr] <= mem_MPORT_479_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_480_en & mem_MPORT_480_mask) begin
      mem[mem_MPORT_480_addr] <= mem_MPORT_480_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_481_en & mem_MPORT_481_mask) begin
      mem[mem_MPORT_481_addr] <= mem_MPORT_481_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_482_en & mem_MPORT_482_mask) begin
      mem[mem_MPORT_482_addr] <= mem_MPORT_482_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_483_en & mem_MPORT_483_mask) begin
      mem[mem_MPORT_483_addr] <= mem_MPORT_483_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_484_en & mem_MPORT_484_mask) begin
      mem[mem_MPORT_484_addr] <= mem_MPORT_484_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_485_en & mem_MPORT_485_mask) begin
      mem[mem_MPORT_485_addr] <= mem_MPORT_485_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_486_en & mem_MPORT_486_mask) begin
      mem[mem_MPORT_486_addr] <= mem_MPORT_486_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_487_en & mem_MPORT_487_mask) begin
      mem[mem_MPORT_487_addr] <= mem_MPORT_487_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_488_en & mem_MPORT_488_mask) begin
      mem[mem_MPORT_488_addr] <= mem_MPORT_488_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_489_en & mem_MPORT_489_mask) begin
      mem[mem_MPORT_489_addr] <= mem_MPORT_489_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_490_en & mem_MPORT_490_mask) begin
      mem[mem_MPORT_490_addr] <= mem_MPORT_490_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_491_en & mem_MPORT_491_mask) begin
      mem[mem_MPORT_491_addr] <= mem_MPORT_491_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_492_en & mem_MPORT_492_mask) begin
      mem[mem_MPORT_492_addr] <= mem_MPORT_492_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_493_en & mem_MPORT_493_mask) begin
      mem[mem_MPORT_493_addr] <= mem_MPORT_493_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_494_en & mem_MPORT_494_mask) begin
      mem[mem_MPORT_494_addr] <= mem_MPORT_494_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_495_en & mem_MPORT_495_mask) begin
      mem[mem_MPORT_495_addr] <= mem_MPORT_495_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_496_en & mem_MPORT_496_mask) begin
      mem[mem_MPORT_496_addr] <= mem_MPORT_496_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_497_en & mem_MPORT_497_mask) begin
      mem[mem_MPORT_497_addr] <= mem_MPORT_497_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_498_en & mem_MPORT_498_mask) begin
      mem[mem_MPORT_498_addr] <= mem_MPORT_498_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_499_en & mem_MPORT_499_mask) begin
      mem[mem_MPORT_499_addr] <= mem_MPORT_499_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_500_en & mem_MPORT_500_mask) begin
      mem[mem_MPORT_500_addr] <= mem_MPORT_500_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_501_en & mem_MPORT_501_mask) begin
      mem[mem_MPORT_501_addr] <= mem_MPORT_501_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_502_en & mem_MPORT_502_mask) begin
      mem[mem_MPORT_502_addr] <= mem_MPORT_502_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_503_en & mem_MPORT_503_mask) begin
      mem[mem_MPORT_503_addr] <= mem_MPORT_503_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_504_en & mem_MPORT_504_mask) begin
      mem[mem_MPORT_504_addr] <= mem_MPORT_504_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_505_en & mem_MPORT_505_mask) begin
      mem[mem_MPORT_505_addr] <= mem_MPORT_505_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_506_en & mem_MPORT_506_mask) begin
      mem[mem_MPORT_506_addr] <= mem_MPORT_506_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_507_en & mem_MPORT_507_mask) begin
      mem[mem_MPORT_507_addr] <= mem_MPORT_507_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_508_en & mem_MPORT_508_mask) begin
      mem[mem_MPORT_508_addr] <= mem_MPORT_508_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_509_en & mem_MPORT_509_mask) begin
      mem[mem_MPORT_509_addr] <= mem_MPORT_509_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_510_en & mem_MPORT_510_mask) begin
      mem[mem_MPORT_510_addr] <= mem_MPORT_510_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_511_en & mem_MPORT_511_mask) begin
      mem[mem_MPORT_511_addr] <= mem_MPORT_511_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_512_en & mem_MPORT_512_mask) begin
      mem[mem_MPORT_512_addr] <= mem_MPORT_512_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_10(
  input         clock,
  input         reset,
  input  [8:0]  io_r_addr,
  output [31:0] io_r_data_0,
  output [31:0] io_r_data_1,
  output [31:0] io_r_data_2,
  output [31:0] io_r_data_3,
  input         io_w_en,
  input  [8:0]  io_w_addr,
  input  [31:0] io_w_data_0,
  input  [31:0] io_w_data_1,
  input  [31:0] io_w_data_2,
  input  [31:0] io_w_data_3,
  input  [3:0]  io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P_80 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P_80 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P_80 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P_80 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
endmodule
module DataBankArray_1(
  input         clock,
  input         reset,
  output        io_read_req_ready,
  input         io_read_req_valid,
  input  [8:0]  io_read_req_bits_set,
  output [31:0] io_read_resp_0_0,
  output [31:0] io_read_resp_0_1,
  output [31:0] io_read_resp_0_2,
  output [31:0] io_read_resp_0_3,
  output [31:0] io_read_resp_1_0,
  output [31:0] io_read_resp_1_1,
  output [31:0] io_read_resp_1_2,
  output [31:0] io_read_resp_1_3,
  output [31:0] io_read_resp_2_0,
  output [31:0] io_read_resp_2_1,
  output [31:0] io_read_resp_2_2,
  output [31:0] io_read_resp_2_3,
  output [31:0] io_read_resp_3_0,
  output [31:0] io_read_resp_3_1,
  output [31:0] io_read_resp_3_2,
  output [31:0] io_read_resp_3_3,
  output        io_write_req_ready,
  input         io_write_req_valid,
  input  [8:0]  io_write_req_bits_set,
  input  [31:0] io_write_req_bits_data_0,
  input  [31:0] io_write_req_bits_data_1,
  input  [31:0] io_write_req_bits_data_2,
  input  [31:0] io_write_req_bits_data_3,
  input  [3:0]  io_write_req_bits_blockMask,
  input  [3:0]  io_write_req_bits_way
);
  wire  dataBanks_0_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_0_reset; // @[SRAM_1.scala 255:31]
  wire [8:0] dataBanks_0_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_0_io_w_en; // @[SRAM_1.scala 255:31]
  wire [8:0] dataBanks_0_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_0_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_reset; // @[SRAM_1.scala 255:31]
  wire [8:0] dataBanks_1_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_io_w_en; // @[SRAM_1.scala 255:31]
  wire [8:0] dataBanks_1_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_1_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_reset; // @[SRAM_1.scala 255:31]
  wire [8:0] dataBanks_2_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_io_w_en; // @[SRAM_1.scala 255:31]
  wire [8:0] dataBanks_2_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_2_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_reset; // @[SRAM_1.scala 255:31]
  wire [8:0] dataBanks_3_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_io_w_en; // @[SRAM_1.scala 255:31]
  wire [8:0] dataBanks_3_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_3_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  ren = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  wire  _wen_T_1 = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  SRAMArray_2P_10 dataBanks_0 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_0_clock),
    .reset(dataBanks_0_reset),
    .io_r_addr(dataBanks_0_io_r_addr),
    .io_r_data_0(dataBanks_0_io_r_data_0),
    .io_r_data_1(dataBanks_0_io_r_data_1),
    .io_r_data_2(dataBanks_0_io_r_data_2),
    .io_r_data_3(dataBanks_0_io_r_data_3),
    .io_w_en(dataBanks_0_io_w_en),
    .io_w_addr(dataBanks_0_io_w_addr),
    .io_w_data_0(dataBanks_0_io_w_data_0),
    .io_w_data_1(dataBanks_0_io_w_data_1),
    .io_w_data_2(dataBanks_0_io_w_data_2),
    .io_w_data_3(dataBanks_0_io_w_data_3),
    .io_w_maskOH(dataBanks_0_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_1 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_1_clock),
    .reset(dataBanks_1_reset),
    .io_r_addr(dataBanks_1_io_r_addr),
    .io_r_data_0(dataBanks_1_io_r_data_0),
    .io_r_data_1(dataBanks_1_io_r_data_1),
    .io_r_data_2(dataBanks_1_io_r_data_2),
    .io_r_data_3(dataBanks_1_io_r_data_3),
    .io_w_en(dataBanks_1_io_w_en),
    .io_w_addr(dataBanks_1_io_w_addr),
    .io_w_data_0(dataBanks_1_io_w_data_0),
    .io_w_data_1(dataBanks_1_io_w_data_1),
    .io_w_data_2(dataBanks_1_io_w_data_2),
    .io_w_data_3(dataBanks_1_io_w_data_3),
    .io_w_maskOH(dataBanks_1_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_2 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_2_clock),
    .reset(dataBanks_2_reset),
    .io_r_addr(dataBanks_2_io_r_addr),
    .io_r_data_0(dataBanks_2_io_r_data_0),
    .io_r_data_1(dataBanks_2_io_r_data_1),
    .io_r_data_2(dataBanks_2_io_r_data_2),
    .io_r_data_3(dataBanks_2_io_r_data_3),
    .io_w_en(dataBanks_2_io_w_en),
    .io_w_addr(dataBanks_2_io_w_addr),
    .io_w_data_0(dataBanks_2_io_w_data_0),
    .io_w_data_1(dataBanks_2_io_w_data_1),
    .io_w_data_2(dataBanks_2_io_w_data_2),
    .io_w_data_3(dataBanks_2_io_w_data_3),
    .io_w_maskOH(dataBanks_2_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_3 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_3_clock),
    .reset(dataBanks_3_reset),
    .io_r_addr(dataBanks_3_io_r_addr),
    .io_r_data_0(dataBanks_3_io_r_data_0),
    .io_r_data_1(dataBanks_3_io_r_data_1),
    .io_r_data_2(dataBanks_3_io_r_data_2),
    .io_r_data_3(dataBanks_3_io_r_data_3),
    .io_w_en(dataBanks_3_io_w_en),
    .io_w_addr(dataBanks_3_io_w_addr),
    .io_w_data_0(dataBanks_3_io_w_data_0),
    .io_w_data_1(dataBanks_3_io_w_data_1),
    .io_w_data_2(dataBanks_3_io_w_data_2),
    .io_w_data_3(dataBanks_3_io_w_data_3),
    .io_w_maskOH(dataBanks_3_io_w_maskOH)
  );
  assign io_read_req_ready = 1'h1; // @[DataBank.scala 46:23]
  assign io_read_resp_0_0 = ren ? dataBanks_0_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_1 = ren ? dataBanks_0_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_2 = ren ? dataBanks_0_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_3 = ren ? dataBanks_0_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_0 = ren ? dataBanks_1_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_1 = ren ? dataBanks_1_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_2 = ren ? dataBanks_1_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_3 = ren ? dataBanks_1_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_0 = ren ? dataBanks_2_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_1 = ren ? dataBanks_2_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_2 = ren ? dataBanks_2_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_3 = ren ? dataBanks_2_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_0 = ren ? dataBanks_3_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_1 = ren ? dataBanks_3_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_2 = ren ? dataBanks_3_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_3 = ren ? dataBanks_3_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_write_req_ready = 1'h1; // @[DataBank.scala 55:28]
  assign dataBanks_0_clock = clock;
  assign dataBanks_0_reset = reset;
  assign dataBanks_0_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_0_io_w_en = io_write_req_bits_way[0] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_0_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_0_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_1_clock = clock;
  assign dataBanks_1_reset = reset;
  assign dataBanks_1_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_1_io_w_en = io_write_req_bits_way[1] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_1_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_1_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_2_clock = clock;
  assign dataBanks_2_reset = reset;
  assign dataBanks_2_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_2_io_w_en = io_write_req_bits_way[2] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_2_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_2_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_3_clock = clock;
  assign dataBanks_3_reset = reset;
  assign dataBanks_3_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_3_io_w_en = io_write_req_bits_way[3] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_3_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_3_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
endmodule
module BankRAM_2P_96(
  input         clock,
  input         reset,
  input  [8:0]  io_r_addr,
  output [18:0] io_r_data,
  input         io_w_en,
  input  [8:0]  io_w_addr,
  input  [18:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [18:0] mem [0:511]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_129_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_130_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_131_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_132_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_133_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_134_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_135_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_136_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_137_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_138_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_139_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_140_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_141_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_142_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_143_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_144_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_145_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_146_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_147_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_148_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_149_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_150_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_151_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_152_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_153_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_154_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_155_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_156_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_157_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_158_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_159_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_160_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_161_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_162_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_163_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_164_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_165_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_166_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_167_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_168_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_169_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_170_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_171_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_172_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_173_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_174_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_175_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_176_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_177_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_178_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_179_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_180_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_181_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_182_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_183_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_184_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_185_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_186_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_187_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_188_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_189_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_190_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_191_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_192_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_193_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_194_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_195_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_196_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_197_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_198_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_199_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_200_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_201_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_202_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_203_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_204_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_205_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_206_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_207_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_208_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_209_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_210_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_211_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_212_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_213_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_214_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_215_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_216_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_217_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_218_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_219_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_220_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_221_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_222_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_223_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_224_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_225_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_226_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_227_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_228_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_229_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_230_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_231_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_232_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_233_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_234_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_235_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_236_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_237_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_238_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_239_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_240_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_241_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_242_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_243_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_244_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_245_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_246_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_247_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_248_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_249_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_250_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_251_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_252_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_253_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_254_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_255_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_256_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_257_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_257_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_257_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_257_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_258_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_258_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_258_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_258_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_259_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_259_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_259_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_259_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_260_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_260_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_260_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_260_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_261_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_261_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_261_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_261_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_262_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_262_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_262_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_262_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_263_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_263_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_263_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_263_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_264_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_264_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_264_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_264_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_265_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_265_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_265_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_265_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_266_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_266_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_266_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_266_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_267_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_267_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_267_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_267_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_268_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_268_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_268_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_268_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_269_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_269_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_269_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_269_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_270_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_270_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_270_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_270_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_271_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_271_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_271_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_271_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_272_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_272_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_272_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_272_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_273_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_273_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_273_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_273_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_274_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_274_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_274_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_274_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_275_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_275_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_275_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_275_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_276_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_276_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_276_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_276_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_277_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_277_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_277_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_277_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_278_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_278_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_278_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_278_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_279_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_279_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_279_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_279_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_280_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_280_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_280_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_280_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_281_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_281_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_281_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_281_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_282_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_282_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_282_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_282_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_283_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_283_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_283_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_283_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_284_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_284_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_284_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_284_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_285_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_285_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_285_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_285_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_286_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_286_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_286_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_286_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_287_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_287_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_287_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_287_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_288_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_288_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_288_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_288_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_289_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_289_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_289_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_289_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_290_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_290_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_290_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_290_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_291_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_291_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_291_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_291_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_292_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_292_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_292_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_292_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_293_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_293_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_293_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_293_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_294_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_294_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_294_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_294_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_295_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_295_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_295_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_295_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_296_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_296_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_296_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_296_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_297_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_297_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_297_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_297_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_298_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_298_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_298_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_298_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_299_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_299_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_299_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_299_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_300_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_300_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_300_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_300_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_301_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_301_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_301_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_301_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_302_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_302_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_302_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_302_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_303_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_303_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_303_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_303_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_304_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_304_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_304_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_304_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_305_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_305_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_305_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_305_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_306_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_306_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_306_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_306_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_307_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_307_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_307_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_307_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_308_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_308_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_308_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_308_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_309_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_309_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_309_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_309_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_310_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_310_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_310_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_310_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_311_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_311_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_311_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_311_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_312_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_312_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_312_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_312_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_313_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_313_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_313_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_313_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_314_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_314_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_314_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_314_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_315_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_315_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_315_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_315_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_316_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_316_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_316_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_316_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_317_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_317_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_317_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_317_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_318_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_318_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_318_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_318_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_319_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_319_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_319_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_319_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_320_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_320_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_320_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_320_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_321_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_321_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_321_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_321_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_322_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_322_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_322_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_322_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_323_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_323_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_323_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_323_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_324_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_324_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_324_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_324_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_325_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_325_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_325_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_325_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_326_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_326_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_326_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_326_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_327_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_327_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_327_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_327_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_328_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_328_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_328_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_328_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_329_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_329_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_329_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_329_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_330_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_330_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_330_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_330_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_331_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_331_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_331_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_331_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_332_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_332_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_332_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_332_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_333_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_333_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_333_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_333_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_334_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_334_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_334_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_334_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_335_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_335_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_335_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_335_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_336_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_336_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_336_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_336_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_337_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_337_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_337_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_337_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_338_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_338_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_338_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_338_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_339_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_339_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_339_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_339_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_340_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_340_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_340_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_340_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_341_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_341_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_341_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_341_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_342_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_342_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_342_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_342_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_343_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_343_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_343_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_343_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_344_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_344_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_344_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_344_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_345_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_345_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_345_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_345_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_346_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_346_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_346_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_346_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_347_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_347_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_347_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_347_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_348_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_348_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_348_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_348_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_349_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_349_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_349_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_349_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_350_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_350_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_350_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_350_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_351_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_351_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_351_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_351_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_352_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_352_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_352_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_352_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_353_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_353_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_353_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_353_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_354_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_354_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_354_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_354_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_355_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_355_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_355_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_355_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_356_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_356_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_356_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_356_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_357_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_357_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_357_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_357_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_358_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_358_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_358_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_358_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_359_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_359_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_359_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_359_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_360_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_360_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_360_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_360_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_361_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_361_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_361_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_361_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_362_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_362_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_362_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_362_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_363_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_363_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_363_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_363_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_364_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_364_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_364_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_364_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_365_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_365_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_365_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_365_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_366_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_366_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_366_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_366_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_367_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_367_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_367_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_367_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_368_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_368_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_368_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_368_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_369_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_369_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_369_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_369_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_370_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_370_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_370_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_370_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_371_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_371_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_371_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_371_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_372_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_372_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_372_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_372_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_373_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_373_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_373_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_373_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_374_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_374_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_374_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_374_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_375_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_375_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_375_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_375_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_376_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_376_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_376_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_376_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_377_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_377_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_377_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_377_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_378_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_378_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_378_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_378_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_379_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_379_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_379_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_379_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_380_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_380_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_380_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_380_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_381_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_381_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_381_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_381_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_382_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_382_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_382_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_382_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_383_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_383_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_383_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_383_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_384_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_384_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_384_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_384_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_385_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_385_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_385_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_385_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_386_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_386_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_386_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_386_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_387_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_387_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_387_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_387_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_388_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_388_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_388_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_388_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_389_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_389_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_389_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_389_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_390_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_390_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_390_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_390_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_391_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_391_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_391_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_391_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_392_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_392_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_392_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_392_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_393_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_393_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_393_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_393_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_394_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_394_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_394_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_394_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_395_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_395_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_395_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_395_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_396_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_396_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_396_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_396_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_397_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_397_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_397_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_397_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_398_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_398_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_398_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_398_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_399_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_399_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_399_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_399_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_400_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_400_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_400_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_400_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_401_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_401_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_401_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_401_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_402_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_402_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_402_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_402_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_403_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_403_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_403_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_403_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_404_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_404_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_404_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_404_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_405_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_405_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_405_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_405_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_406_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_406_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_406_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_406_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_407_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_407_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_407_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_407_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_408_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_408_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_408_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_408_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_409_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_409_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_409_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_409_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_410_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_410_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_410_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_410_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_411_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_411_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_411_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_411_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_412_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_412_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_412_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_412_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_413_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_413_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_413_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_413_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_414_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_414_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_414_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_414_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_415_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_415_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_415_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_415_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_416_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_416_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_416_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_416_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_417_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_417_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_417_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_417_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_418_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_418_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_418_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_418_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_419_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_419_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_419_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_419_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_420_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_420_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_420_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_420_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_421_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_421_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_421_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_421_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_422_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_422_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_422_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_422_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_423_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_423_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_423_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_423_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_424_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_424_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_424_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_424_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_425_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_425_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_425_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_425_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_426_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_426_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_426_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_426_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_427_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_427_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_427_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_427_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_428_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_428_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_428_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_428_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_429_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_429_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_429_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_429_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_430_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_430_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_430_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_430_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_431_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_431_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_431_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_431_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_432_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_432_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_432_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_432_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_433_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_433_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_433_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_433_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_434_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_434_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_434_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_434_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_435_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_435_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_435_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_435_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_436_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_436_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_436_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_436_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_437_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_437_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_437_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_437_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_438_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_438_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_438_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_438_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_439_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_439_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_439_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_439_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_440_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_440_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_440_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_440_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_441_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_441_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_441_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_441_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_442_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_442_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_442_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_442_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_443_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_443_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_443_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_443_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_444_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_444_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_444_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_444_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_445_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_445_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_445_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_445_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_446_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_446_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_446_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_446_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_447_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_447_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_447_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_447_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_448_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_448_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_448_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_448_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_449_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_449_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_449_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_449_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_450_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_450_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_450_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_450_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_451_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_451_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_451_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_451_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_452_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_452_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_452_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_452_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_453_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_453_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_453_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_453_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_454_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_454_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_454_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_454_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_455_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_455_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_455_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_455_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_456_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_456_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_456_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_456_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_457_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_457_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_457_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_457_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_458_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_458_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_458_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_458_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_459_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_459_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_459_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_459_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_460_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_460_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_460_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_460_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_461_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_461_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_461_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_461_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_462_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_462_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_462_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_462_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_463_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_463_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_463_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_463_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_464_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_464_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_464_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_464_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_465_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_465_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_465_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_465_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_466_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_466_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_466_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_466_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_467_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_467_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_467_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_467_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_468_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_468_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_468_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_468_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_469_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_469_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_469_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_469_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_470_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_470_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_470_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_470_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_471_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_471_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_471_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_471_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_472_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_472_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_472_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_472_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_473_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_473_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_473_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_473_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_474_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_474_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_474_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_474_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_475_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_475_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_475_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_475_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_476_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_476_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_476_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_476_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_477_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_477_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_477_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_477_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_478_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_478_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_478_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_478_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_479_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_479_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_479_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_479_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_480_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_480_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_480_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_480_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_481_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_481_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_481_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_481_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_482_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_482_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_482_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_482_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_483_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_483_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_483_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_483_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_484_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_484_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_484_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_484_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_485_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_485_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_485_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_485_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_486_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_486_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_486_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_486_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_487_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_487_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_487_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_487_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_488_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_488_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_488_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_488_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_489_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_489_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_489_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_489_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_490_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_490_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_490_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_490_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_491_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_491_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_491_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_491_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_492_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_492_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_492_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_492_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_493_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_493_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_493_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_493_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_494_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_494_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_494_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_494_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_495_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_495_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_495_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_495_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_496_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_496_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_496_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_496_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_497_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_497_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_497_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_497_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_498_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_498_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_498_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_498_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_499_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_499_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_499_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_499_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_500_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_500_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_500_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_500_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_501_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_501_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_501_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_501_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_502_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_502_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_502_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_502_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_503_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_503_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_503_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_503_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_504_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_504_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_504_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_504_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_505_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_505_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_505_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_505_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_506_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_506_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_506_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_506_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_507_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_507_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_507_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_507_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_508_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_508_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_508_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_508_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_509_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_509_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_509_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_509_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_510_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_510_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_510_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_510_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_511_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_511_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_511_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_511_en; // @[SRAM_1.scala 63:26]
  wire [18:0] mem_MPORT_512_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_512_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_512_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_512_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [8:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 19'h0;
  assign mem_MPORT_addr = 9'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 19'h0;
  assign mem_MPORT_1_addr = 9'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 19'h0;
  assign mem_MPORT_2_addr = 9'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 19'h0;
  assign mem_MPORT_3_addr = 9'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 19'h0;
  assign mem_MPORT_4_addr = 9'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 19'h0;
  assign mem_MPORT_5_addr = 9'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 19'h0;
  assign mem_MPORT_6_addr = 9'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 19'h0;
  assign mem_MPORT_7_addr = 9'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 19'h0;
  assign mem_MPORT_8_addr = 9'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 19'h0;
  assign mem_MPORT_9_addr = 9'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 19'h0;
  assign mem_MPORT_10_addr = 9'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 19'h0;
  assign mem_MPORT_11_addr = 9'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 19'h0;
  assign mem_MPORT_12_addr = 9'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 19'h0;
  assign mem_MPORT_13_addr = 9'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 19'h0;
  assign mem_MPORT_14_addr = 9'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 19'h0;
  assign mem_MPORT_15_addr = 9'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 19'h0;
  assign mem_MPORT_16_addr = 9'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 19'h0;
  assign mem_MPORT_17_addr = 9'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 19'h0;
  assign mem_MPORT_18_addr = 9'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 19'h0;
  assign mem_MPORT_19_addr = 9'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 19'h0;
  assign mem_MPORT_20_addr = 9'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 19'h0;
  assign mem_MPORT_21_addr = 9'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 19'h0;
  assign mem_MPORT_22_addr = 9'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 19'h0;
  assign mem_MPORT_23_addr = 9'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 19'h0;
  assign mem_MPORT_24_addr = 9'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 19'h0;
  assign mem_MPORT_25_addr = 9'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 19'h0;
  assign mem_MPORT_26_addr = 9'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 19'h0;
  assign mem_MPORT_27_addr = 9'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 19'h0;
  assign mem_MPORT_28_addr = 9'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 19'h0;
  assign mem_MPORT_29_addr = 9'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 19'h0;
  assign mem_MPORT_30_addr = 9'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 19'h0;
  assign mem_MPORT_31_addr = 9'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 19'h0;
  assign mem_MPORT_32_addr = 9'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 19'h0;
  assign mem_MPORT_33_addr = 9'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 19'h0;
  assign mem_MPORT_34_addr = 9'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 19'h0;
  assign mem_MPORT_35_addr = 9'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 19'h0;
  assign mem_MPORT_36_addr = 9'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 19'h0;
  assign mem_MPORT_37_addr = 9'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 19'h0;
  assign mem_MPORT_38_addr = 9'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 19'h0;
  assign mem_MPORT_39_addr = 9'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 19'h0;
  assign mem_MPORT_40_addr = 9'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 19'h0;
  assign mem_MPORT_41_addr = 9'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 19'h0;
  assign mem_MPORT_42_addr = 9'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 19'h0;
  assign mem_MPORT_43_addr = 9'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 19'h0;
  assign mem_MPORT_44_addr = 9'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 19'h0;
  assign mem_MPORT_45_addr = 9'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 19'h0;
  assign mem_MPORT_46_addr = 9'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 19'h0;
  assign mem_MPORT_47_addr = 9'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 19'h0;
  assign mem_MPORT_48_addr = 9'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 19'h0;
  assign mem_MPORT_49_addr = 9'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 19'h0;
  assign mem_MPORT_50_addr = 9'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 19'h0;
  assign mem_MPORT_51_addr = 9'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 19'h0;
  assign mem_MPORT_52_addr = 9'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 19'h0;
  assign mem_MPORT_53_addr = 9'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 19'h0;
  assign mem_MPORT_54_addr = 9'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 19'h0;
  assign mem_MPORT_55_addr = 9'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 19'h0;
  assign mem_MPORT_56_addr = 9'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 19'h0;
  assign mem_MPORT_57_addr = 9'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 19'h0;
  assign mem_MPORT_58_addr = 9'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 19'h0;
  assign mem_MPORT_59_addr = 9'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 19'h0;
  assign mem_MPORT_60_addr = 9'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 19'h0;
  assign mem_MPORT_61_addr = 9'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 19'h0;
  assign mem_MPORT_62_addr = 9'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 19'h0;
  assign mem_MPORT_63_addr = 9'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 19'h0;
  assign mem_MPORT_64_addr = 9'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 19'h0;
  assign mem_MPORT_65_addr = 9'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 19'h0;
  assign mem_MPORT_66_addr = 9'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 19'h0;
  assign mem_MPORT_67_addr = 9'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 19'h0;
  assign mem_MPORT_68_addr = 9'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 19'h0;
  assign mem_MPORT_69_addr = 9'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 19'h0;
  assign mem_MPORT_70_addr = 9'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 19'h0;
  assign mem_MPORT_71_addr = 9'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 19'h0;
  assign mem_MPORT_72_addr = 9'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 19'h0;
  assign mem_MPORT_73_addr = 9'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 19'h0;
  assign mem_MPORT_74_addr = 9'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 19'h0;
  assign mem_MPORT_75_addr = 9'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 19'h0;
  assign mem_MPORT_76_addr = 9'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 19'h0;
  assign mem_MPORT_77_addr = 9'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 19'h0;
  assign mem_MPORT_78_addr = 9'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 19'h0;
  assign mem_MPORT_79_addr = 9'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 19'h0;
  assign mem_MPORT_80_addr = 9'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 19'h0;
  assign mem_MPORT_81_addr = 9'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 19'h0;
  assign mem_MPORT_82_addr = 9'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 19'h0;
  assign mem_MPORT_83_addr = 9'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 19'h0;
  assign mem_MPORT_84_addr = 9'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 19'h0;
  assign mem_MPORT_85_addr = 9'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 19'h0;
  assign mem_MPORT_86_addr = 9'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 19'h0;
  assign mem_MPORT_87_addr = 9'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 19'h0;
  assign mem_MPORT_88_addr = 9'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 19'h0;
  assign mem_MPORT_89_addr = 9'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 19'h0;
  assign mem_MPORT_90_addr = 9'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 19'h0;
  assign mem_MPORT_91_addr = 9'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 19'h0;
  assign mem_MPORT_92_addr = 9'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 19'h0;
  assign mem_MPORT_93_addr = 9'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 19'h0;
  assign mem_MPORT_94_addr = 9'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 19'h0;
  assign mem_MPORT_95_addr = 9'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 19'h0;
  assign mem_MPORT_96_addr = 9'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 19'h0;
  assign mem_MPORT_97_addr = 9'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 19'h0;
  assign mem_MPORT_98_addr = 9'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 19'h0;
  assign mem_MPORT_99_addr = 9'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 19'h0;
  assign mem_MPORT_100_addr = 9'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 19'h0;
  assign mem_MPORT_101_addr = 9'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 19'h0;
  assign mem_MPORT_102_addr = 9'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 19'h0;
  assign mem_MPORT_103_addr = 9'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 19'h0;
  assign mem_MPORT_104_addr = 9'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 19'h0;
  assign mem_MPORT_105_addr = 9'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 19'h0;
  assign mem_MPORT_106_addr = 9'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 19'h0;
  assign mem_MPORT_107_addr = 9'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 19'h0;
  assign mem_MPORT_108_addr = 9'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 19'h0;
  assign mem_MPORT_109_addr = 9'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 19'h0;
  assign mem_MPORT_110_addr = 9'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 19'h0;
  assign mem_MPORT_111_addr = 9'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 19'h0;
  assign mem_MPORT_112_addr = 9'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 19'h0;
  assign mem_MPORT_113_addr = 9'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 19'h0;
  assign mem_MPORT_114_addr = 9'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 19'h0;
  assign mem_MPORT_115_addr = 9'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 19'h0;
  assign mem_MPORT_116_addr = 9'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 19'h0;
  assign mem_MPORT_117_addr = 9'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 19'h0;
  assign mem_MPORT_118_addr = 9'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 19'h0;
  assign mem_MPORT_119_addr = 9'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 19'h0;
  assign mem_MPORT_120_addr = 9'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 19'h0;
  assign mem_MPORT_121_addr = 9'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 19'h0;
  assign mem_MPORT_122_addr = 9'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 19'h0;
  assign mem_MPORT_123_addr = 9'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 19'h0;
  assign mem_MPORT_124_addr = 9'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 19'h0;
  assign mem_MPORT_125_addr = 9'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 19'h0;
  assign mem_MPORT_126_addr = 9'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 19'h0;
  assign mem_MPORT_127_addr = 9'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 19'h0;
  assign mem_MPORT_128_addr = 9'h80;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = reset;
  assign mem_MPORT_129_data = 19'h0;
  assign mem_MPORT_129_addr = 9'h81;
  assign mem_MPORT_129_mask = 1'h1;
  assign mem_MPORT_129_en = reset;
  assign mem_MPORT_130_data = 19'h0;
  assign mem_MPORT_130_addr = 9'h82;
  assign mem_MPORT_130_mask = 1'h1;
  assign mem_MPORT_130_en = reset;
  assign mem_MPORT_131_data = 19'h0;
  assign mem_MPORT_131_addr = 9'h83;
  assign mem_MPORT_131_mask = 1'h1;
  assign mem_MPORT_131_en = reset;
  assign mem_MPORT_132_data = 19'h0;
  assign mem_MPORT_132_addr = 9'h84;
  assign mem_MPORT_132_mask = 1'h1;
  assign mem_MPORT_132_en = reset;
  assign mem_MPORT_133_data = 19'h0;
  assign mem_MPORT_133_addr = 9'h85;
  assign mem_MPORT_133_mask = 1'h1;
  assign mem_MPORT_133_en = reset;
  assign mem_MPORT_134_data = 19'h0;
  assign mem_MPORT_134_addr = 9'h86;
  assign mem_MPORT_134_mask = 1'h1;
  assign mem_MPORT_134_en = reset;
  assign mem_MPORT_135_data = 19'h0;
  assign mem_MPORT_135_addr = 9'h87;
  assign mem_MPORT_135_mask = 1'h1;
  assign mem_MPORT_135_en = reset;
  assign mem_MPORT_136_data = 19'h0;
  assign mem_MPORT_136_addr = 9'h88;
  assign mem_MPORT_136_mask = 1'h1;
  assign mem_MPORT_136_en = reset;
  assign mem_MPORT_137_data = 19'h0;
  assign mem_MPORT_137_addr = 9'h89;
  assign mem_MPORT_137_mask = 1'h1;
  assign mem_MPORT_137_en = reset;
  assign mem_MPORT_138_data = 19'h0;
  assign mem_MPORT_138_addr = 9'h8a;
  assign mem_MPORT_138_mask = 1'h1;
  assign mem_MPORT_138_en = reset;
  assign mem_MPORT_139_data = 19'h0;
  assign mem_MPORT_139_addr = 9'h8b;
  assign mem_MPORT_139_mask = 1'h1;
  assign mem_MPORT_139_en = reset;
  assign mem_MPORT_140_data = 19'h0;
  assign mem_MPORT_140_addr = 9'h8c;
  assign mem_MPORT_140_mask = 1'h1;
  assign mem_MPORT_140_en = reset;
  assign mem_MPORT_141_data = 19'h0;
  assign mem_MPORT_141_addr = 9'h8d;
  assign mem_MPORT_141_mask = 1'h1;
  assign mem_MPORT_141_en = reset;
  assign mem_MPORT_142_data = 19'h0;
  assign mem_MPORT_142_addr = 9'h8e;
  assign mem_MPORT_142_mask = 1'h1;
  assign mem_MPORT_142_en = reset;
  assign mem_MPORT_143_data = 19'h0;
  assign mem_MPORT_143_addr = 9'h8f;
  assign mem_MPORT_143_mask = 1'h1;
  assign mem_MPORT_143_en = reset;
  assign mem_MPORT_144_data = 19'h0;
  assign mem_MPORT_144_addr = 9'h90;
  assign mem_MPORT_144_mask = 1'h1;
  assign mem_MPORT_144_en = reset;
  assign mem_MPORT_145_data = 19'h0;
  assign mem_MPORT_145_addr = 9'h91;
  assign mem_MPORT_145_mask = 1'h1;
  assign mem_MPORT_145_en = reset;
  assign mem_MPORT_146_data = 19'h0;
  assign mem_MPORT_146_addr = 9'h92;
  assign mem_MPORT_146_mask = 1'h1;
  assign mem_MPORT_146_en = reset;
  assign mem_MPORT_147_data = 19'h0;
  assign mem_MPORT_147_addr = 9'h93;
  assign mem_MPORT_147_mask = 1'h1;
  assign mem_MPORT_147_en = reset;
  assign mem_MPORT_148_data = 19'h0;
  assign mem_MPORT_148_addr = 9'h94;
  assign mem_MPORT_148_mask = 1'h1;
  assign mem_MPORT_148_en = reset;
  assign mem_MPORT_149_data = 19'h0;
  assign mem_MPORT_149_addr = 9'h95;
  assign mem_MPORT_149_mask = 1'h1;
  assign mem_MPORT_149_en = reset;
  assign mem_MPORT_150_data = 19'h0;
  assign mem_MPORT_150_addr = 9'h96;
  assign mem_MPORT_150_mask = 1'h1;
  assign mem_MPORT_150_en = reset;
  assign mem_MPORT_151_data = 19'h0;
  assign mem_MPORT_151_addr = 9'h97;
  assign mem_MPORT_151_mask = 1'h1;
  assign mem_MPORT_151_en = reset;
  assign mem_MPORT_152_data = 19'h0;
  assign mem_MPORT_152_addr = 9'h98;
  assign mem_MPORT_152_mask = 1'h1;
  assign mem_MPORT_152_en = reset;
  assign mem_MPORT_153_data = 19'h0;
  assign mem_MPORT_153_addr = 9'h99;
  assign mem_MPORT_153_mask = 1'h1;
  assign mem_MPORT_153_en = reset;
  assign mem_MPORT_154_data = 19'h0;
  assign mem_MPORT_154_addr = 9'h9a;
  assign mem_MPORT_154_mask = 1'h1;
  assign mem_MPORT_154_en = reset;
  assign mem_MPORT_155_data = 19'h0;
  assign mem_MPORT_155_addr = 9'h9b;
  assign mem_MPORT_155_mask = 1'h1;
  assign mem_MPORT_155_en = reset;
  assign mem_MPORT_156_data = 19'h0;
  assign mem_MPORT_156_addr = 9'h9c;
  assign mem_MPORT_156_mask = 1'h1;
  assign mem_MPORT_156_en = reset;
  assign mem_MPORT_157_data = 19'h0;
  assign mem_MPORT_157_addr = 9'h9d;
  assign mem_MPORT_157_mask = 1'h1;
  assign mem_MPORT_157_en = reset;
  assign mem_MPORT_158_data = 19'h0;
  assign mem_MPORT_158_addr = 9'h9e;
  assign mem_MPORT_158_mask = 1'h1;
  assign mem_MPORT_158_en = reset;
  assign mem_MPORT_159_data = 19'h0;
  assign mem_MPORT_159_addr = 9'h9f;
  assign mem_MPORT_159_mask = 1'h1;
  assign mem_MPORT_159_en = reset;
  assign mem_MPORT_160_data = 19'h0;
  assign mem_MPORT_160_addr = 9'ha0;
  assign mem_MPORT_160_mask = 1'h1;
  assign mem_MPORT_160_en = reset;
  assign mem_MPORT_161_data = 19'h0;
  assign mem_MPORT_161_addr = 9'ha1;
  assign mem_MPORT_161_mask = 1'h1;
  assign mem_MPORT_161_en = reset;
  assign mem_MPORT_162_data = 19'h0;
  assign mem_MPORT_162_addr = 9'ha2;
  assign mem_MPORT_162_mask = 1'h1;
  assign mem_MPORT_162_en = reset;
  assign mem_MPORT_163_data = 19'h0;
  assign mem_MPORT_163_addr = 9'ha3;
  assign mem_MPORT_163_mask = 1'h1;
  assign mem_MPORT_163_en = reset;
  assign mem_MPORT_164_data = 19'h0;
  assign mem_MPORT_164_addr = 9'ha4;
  assign mem_MPORT_164_mask = 1'h1;
  assign mem_MPORT_164_en = reset;
  assign mem_MPORT_165_data = 19'h0;
  assign mem_MPORT_165_addr = 9'ha5;
  assign mem_MPORT_165_mask = 1'h1;
  assign mem_MPORT_165_en = reset;
  assign mem_MPORT_166_data = 19'h0;
  assign mem_MPORT_166_addr = 9'ha6;
  assign mem_MPORT_166_mask = 1'h1;
  assign mem_MPORT_166_en = reset;
  assign mem_MPORT_167_data = 19'h0;
  assign mem_MPORT_167_addr = 9'ha7;
  assign mem_MPORT_167_mask = 1'h1;
  assign mem_MPORT_167_en = reset;
  assign mem_MPORT_168_data = 19'h0;
  assign mem_MPORT_168_addr = 9'ha8;
  assign mem_MPORT_168_mask = 1'h1;
  assign mem_MPORT_168_en = reset;
  assign mem_MPORT_169_data = 19'h0;
  assign mem_MPORT_169_addr = 9'ha9;
  assign mem_MPORT_169_mask = 1'h1;
  assign mem_MPORT_169_en = reset;
  assign mem_MPORT_170_data = 19'h0;
  assign mem_MPORT_170_addr = 9'haa;
  assign mem_MPORT_170_mask = 1'h1;
  assign mem_MPORT_170_en = reset;
  assign mem_MPORT_171_data = 19'h0;
  assign mem_MPORT_171_addr = 9'hab;
  assign mem_MPORT_171_mask = 1'h1;
  assign mem_MPORT_171_en = reset;
  assign mem_MPORT_172_data = 19'h0;
  assign mem_MPORT_172_addr = 9'hac;
  assign mem_MPORT_172_mask = 1'h1;
  assign mem_MPORT_172_en = reset;
  assign mem_MPORT_173_data = 19'h0;
  assign mem_MPORT_173_addr = 9'had;
  assign mem_MPORT_173_mask = 1'h1;
  assign mem_MPORT_173_en = reset;
  assign mem_MPORT_174_data = 19'h0;
  assign mem_MPORT_174_addr = 9'hae;
  assign mem_MPORT_174_mask = 1'h1;
  assign mem_MPORT_174_en = reset;
  assign mem_MPORT_175_data = 19'h0;
  assign mem_MPORT_175_addr = 9'haf;
  assign mem_MPORT_175_mask = 1'h1;
  assign mem_MPORT_175_en = reset;
  assign mem_MPORT_176_data = 19'h0;
  assign mem_MPORT_176_addr = 9'hb0;
  assign mem_MPORT_176_mask = 1'h1;
  assign mem_MPORT_176_en = reset;
  assign mem_MPORT_177_data = 19'h0;
  assign mem_MPORT_177_addr = 9'hb1;
  assign mem_MPORT_177_mask = 1'h1;
  assign mem_MPORT_177_en = reset;
  assign mem_MPORT_178_data = 19'h0;
  assign mem_MPORT_178_addr = 9'hb2;
  assign mem_MPORT_178_mask = 1'h1;
  assign mem_MPORT_178_en = reset;
  assign mem_MPORT_179_data = 19'h0;
  assign mem_MPORT_179_addr = 9'hb3;
  assign mem_MPORT_179_mask = 1'h1;
  assign mem_MPORT_179_en = reset;
  assign mem_MPORT_180_data = 19'h0;
  assign mem_MPORT_180_addr = 9'hb4;
  assign mem_MPORT_180_mask = 1'h1;
  assign mem_MPORT_180_en = reset;
  assign mem_MPORT_181_data = 19'h0;
  assign mem_MPORT_181_addr = 9'hb5;
  assign mem_MPORT_181_mask = 1'h1;
  assign mem_MPORT_181_en = reset;
  assign mem_MPORT_182_data = 19'h0;
  assign mem_MPORT_182_addr = 9'hb6;
  assign mem_MPORT_182_mask = 1'h1;
  assign mem_MPORT_182_en = reset;
  assign mem_MPORT_183_data = 19'h0;
  assign mem_MPORT_183_addr = 9'hb7;
  assign mem_MPORT_183_mask = 1'h1;
  assign mem_MPORT_183_en = reset;
  assign mem_MPORT_184_data = 19'h0;
  assign mem_MPORT_184_addr = 9'hb8;
  assign mem_MPORT_184_mask = 1'h1;
  assign mem_MPORT_184_en = reset;
  assign mem_MPORT_185_data = 19'h0;
  assign mem_MPORT_185_addr = 9'hb9;
  assign mem_MPORT_185_mask = 1'h1;
  assign mem_MPORT_185_en = reset;
  assign mem_MPORT_186_data = 19'h0;
  assign mem_MPORT_186_addr = 9'hba;
  assign mem_MPORT_186_mask = 1'h1;
  assign mem_MPORT_186_en = reset;
  assign mem_MPORT_187_data = 19'h0;
  assign mem_MPORT_187_addr = 9'hbb;
  assign mem_MPORT_187_mask = 1'h1;
  assign mem_MPORT_187_en = reset;
  assign mem_MPORT_188_data = 19'h0;
  assign mem_MPORT_188_addr = 9'hbc;
  assign mem_MPORT_188_mask = 1'h1;
  assign mem_MPORT_188_en = reset;
  assign mem_MPORT_189_data = 19'h0;
  assign mem_MPORT_189_addr = 9'hbd;
  assign mem_MPORT_189_mask = 1'h1;
  assign mem_MPORT_189_en = reset;
  assign mem_MPORT_190_data = 19'h0;
  assign mem_MPORT_190_addr = 9'hbe;
  assign mem_MPORT_190_mask = 1'h1;
  assign mem_MPORT_190_en = reset;
  assign mem_MPORT_191_data = 19'h0;
  assign mem_MPORT_191_addr = 9'hbf;
  assign mem_MPORT_191_mask = 1'h1;
  assign mem_MPORT_191_en = reset;
  assign mem_MPORT_192_data = 19'h0;
  assign mem_MPORT_192_addr = 9'hc0;
  assign mem_MPORT_192_mask = 1'h1;
  assign mem_MPORT_192_en = reset;
  assign mem_MPORT_193_data = 19'h0;
  assign mem_MPORT_193_addr = 9'hc1;
  assign mem_MPORT_193_mask = 1'h1;
  assign mem_MPORT_193_en = reset;
  assign mem_MPORT_194_data = 19'h0;
  assign mem_MPORT_194_addr = 9'hc2;
  assign mem_MPORT_194_mask = 1'h1;
  assign mem_MPORT_194_en = reset;
  assign mem_MPORT_195_data = 19'h0;
  assign mem_MPORT_195_addr = 9'hc3;
  assign mem_MPORT_195_mask = 1'h1;
  assign mem_MPORT_195_en = reset;
  assign mem_MPORT_196_data = 19'h0;
  assign mem_MPORT_196_addr = 9'hc4;
  assign mem_MPORT_196_mask = 1'h1;
  assign mem_MPORT_196_en = reset;
  assign mem_MPORT_197_data = 19'h0;
  assign mem_MPORT_197_addr = 9'hc5;
  assign mem_MPORT_197_mask = 1'h1;
  assign mem_MPORT_197_en = reset;
  assign mem_MPORT_198_data = 19'h0;
  assign mem_MPORT_198_addr = 9'hc6;
  assign mem_MPORT_198_mask = 1'h1;
  assign mem_MPORT_198_en = reset;
  assign mem_MPORT_199_data = 19'h0;
  assign mem_MPORT_199_addr = 9'hc7;
  assign mem_MPORT_199_mask = 1'h1;
  assign mem_MPORT_199_en = reset;
  assign mem_MPORT_200_data = 19'h0;
  assign mem_MPORT_200_addr = 9'hc8;
  assign mem_MPORT_200_mask = 1'h1;
  assign mem_MPORT_200_en = reset;
  assign mem_MPORT_201_data = 19'h0;
  assign mem_MPORT_201_addr = 9'hc9;
  assign mem_MPORT_201_mask = 1'h1;
  assign mem_MPORT_201_en = reset;
  assign mem_MPORT_202_data = 19'h0;
  assign mem_MPORT_202_addr = 9'hca;
  assign mem_MPORT_202_mask = 1'h1;
  assign mem_MPORT_202_en = reset;
  assign mem_MPORT_203_data = 19'h0;
  assign mem_MPORT_203_addr = 9'hcb;
  assign mem_MPORT_203_mask = 1'h1;
  assign mem_MPORT_203_en = reset;
  assign mem_MPORT_204_data = 19'h0;
  assign mem_MPORT_204_addr = 9'hcc;
  assign mem_MPORT_204_mask = 1'h1;
  assign mem_MPORT_204_en = reset;
  assign mem_MPORT_205_data = 19'h0;
  assign mem_MPORT_205_addr = 9'hcd;
  assign mem_MPORT_205_mask = 1'h1;
  assign mem_MPORT_205_en = reset;
  assign mem_MPORT_206_data = 19'h0;
  assign mem_MPORT_206_addr = 9'hce;
  assign mem_MPORT_206_mask = 1'h1;
  assign mem_MPORT_206_en = reset;
  assign mem_MPORT_207_data = 19'h0;
  assign mem_MPORT_207_addr = 9'hcf;
  assign mem_MPORT_207_mask = 1'h1;
  assign mem_MPORT_207_en = reset;
  assign mem_MPORT_208_data = 19'h0;
  assign mem_MPORT_208_addr = 9'hd0;
  assign mem_MPORT_208_mask = 1'h1;
  assign mem_MPORT_208_en = reset;
  assign mem_MPORT_209_data = 19'h0;
  assign mem_MPORT_209_addr = 9'hd1;
  assign mem_MPORT_209_mask = 1'h1;
  assign mem_MPORT_209_en = reset;
  assign mem_MPORT_210_data = 19'h0;
  assign mem_MPORT_210_addr = 9'hd2;
  assign mem_MPORT_210_mask = 1'h1;
  assign mem_MPORT_210_en = reset;
  assign mem_MPORT_211_data = 19'h0;
  assign mem_MPORT_211_addr = 9'hd3;
  assign mem_MPORT_211_mask = 1'h1;
  assign mem_MPORT_211_en = reset;
  assign mem_MPORT_212_data = 19'h0;
  assign mem_MPORT_212_addr = 9'hd4;
  assign mem_MPORT_212_mask = 1'h1;
  assign mem_MPORT_212_en = reset;
  assign mem_MPORT_213_data = 19'h0;
  assign mem_MPORT_213_addr = 9'hd5;
  assign mem_MPORT_213_mask = 1'h1;
  assign mem_MPORT_213_en = reset;
  assign mem_MPORT_214_data = 19'h0;
  assign mem_MPORT_214_addr = 9'hd6;
  assign mem_MPORT_214_mask = 1'h1;
  assign mem_MPORT_214_en = reset;
  assign mem_MPORT_215_data = 19'h0;
  assign mem_MPORT_215_addr = 9'hd7;
  assign mem_MPORT_215_mask = 1'h1;
  assign mem_MPORT_215_en = reset;
  assign mem_MPORT_216_data = 19'h0;
  assign mem_MPORT_216_addr = 9'hd8;
  assign mem_MPORT_216_mask = 1'h1;
  assign mem_MPORT_216_en = reset;
  assign mem_MPORT_217_data = 19'h0;
  assign mem_MPORT_217_addr = 9'hd9;
  assign mem_MPORT_217_mask = 1'h1;
  assign mem_MPORT_217_en = reset;
  assign mem_MPORT_218_data = 19'h0;
  assign mem_MPORT_218_addr = 9'hda;
  assign mem_MPORT_218_mask = 1'h1;
  assign mem_MPORT_218_en = reset;
  assign mem_MPORT_219_data = 19'h0;
  assign mem_MPORT_219_addr = 9'hdb;
  assign mem_MPORT_219_mask = 1'h1;
  assign mem_MPORT_219_en = reset;
  assign mem_MPORT_220_data = 19'h0;
  assign mem_MPORT_220_addr = 9'hdc;
  assign mem_MPORT_220_mask = 1'h1;
  assign mem_MPORT_220_en = reset;
  assign mem_MPORT_221_data = 19'h0;
  assign mem_MPORT_221_addr = 9'hdd;
  assign mem_MPORT_221_mask = 1'h1;
  assign mem_MPORT_221_en = reset;
  assign mem_MPORT_222_data = 19'h0;
  assign mem_MPORT_222_addr = 9'hde;
  assign mem_MPORT_222_mask = 1'h1;
  assign mem_MPORT_222_en = reset;
  assign mem_MPORT_223_data = 19'h0;
  assign mem_MPORT_223_addr = 9'hdf;
  assign mem_MPORT_223_mask = 1'h1;
  assign mem_MPORT_223_en = reset;
  assign mem_MPORT_224_data = 19'h0;
  assign mem_MPORT_224_addr = 9'he0;
  assign mem_MPORT_224_mask = 1'h1;
  assign mem_MPORT_224_en = reset;
  assign mem_MPORT_225_data = 19'h0;
  assign mem_MPORT_225_addr = 9'he1;
  assign mem_MPORT_225_mask = 1'h1;
  assign mem_MPORT_225_en = reset;
  assign mem_MPORT_226_data = 19'h0;
  assign mem_MPORT_226_addr = 9'he2;
  assign mem_MPORT_226_mask = 1'h1;
  assign mem_MPORT_226_en = reset;
  assign mem_MPORT_227_data = 19'h0;
  assign mem_MPORT_227_addr = 9'he3;
  assign mem_MPORT_227_mask = 1'h1;
  assign mem_MPORT_227_en = reset;
  assign mem_MPORT_228_data = 19'h0;
  assign mem_MPORT_228_addr = 9'he4;
  assign mem_MPORT_228_mask = 1'h1;
  assign mem_MPORT_228_en = reset;
  assign mem_MPORT_229_data = 19'h0;
  assign mem_MPORT_229_addr = 9'he5;
  assign mem_MPORT_229_mask = 1'h1;
  assign mem_MPORT_229_en = reset;
  assign mem_MPORT_230_data = 19'h0;
  assign mem_MPORT_230_addr = 9'he6;
  assign mem_MPORT_230_mask = 1'h1;
  assign mem_MPORT_230_en = reset;
  assign mem_MPORT_231_data = 19'h0;
  assign mem_MPORT_231_addr = 9'he7;
  assign mem_MPORT_231_mask = 1'h1;
  assign mem_MPORT_231_en = reset;
  assign mem_MPORT_232_data = 19'h0;
  assign mem_MPORT_232_addr = 9'he8;
  assign mem_MPORT_232_mask = 1'h1;
  assign mem_MPORT_232_en = reset;
  assign mem_MPORT_233_data = 19'h0;
  assign mem_MPORT_233_addr = 9'he9;
  assign mem_MPORT_233_mask = 1'h1;
  assign mem_MPORT_233_en = reset;
  assign mem_MPORT_234_data = 19'h0;
  assign mem_MPORT_234_addr = 9'hea;
  assign mem_MPORT_234_mask = 1'h1;
  assign mem_MPORT_234_en = reset;
  assign mem_MPORT_235_data = 19'h0;
  assign mem_MPORT_235_addr = 9'heb;
  assign mem_MPORT_235_mask = 1'h1;
  assign mem_MPORT_235_en = reset;
  assign mem_MPORT_236_data = 19'h0;
  assign mem_MPORT_236_addr = 9'hec;
  assign mem_MPORT_236_mask = 1'h1;
  assign mem_MPORT_236_en = reset;
  assign mem_MPORT_237_data = 19'h0;
  assign mem_MPORT_237_addr = 9'hed;
  assign mem_MPORT_237_mask = 1'h1;
  assign mem_MPORT_237_en = reset;
  assign mem_MPORT_238_data = 19'h0;
  assign mem_MPORT_238_addr = 9'hee;
  assign mem_MPORT_238_mask = 1'h1;
  assign mem_MPORT_238_en = reset;
  assign mem_MPORT_239_data = 19'h0;
  assign mem_MPORT_239_addr = 9'hef;
  assign mem_MPORT_239_mask = 1'h1;
  assign mem_MPORT_239_en = reset;
  assign mem_MPORT_240_data = 19'h0;
  assign mem_MPORT_240_addr = 9'hf0;
  assign mem_MPORT_240_mask = 1'h1;
  assign mem_MPORT_240_en = reset;
  assign mem_MPORT_241_data = 19'h0;
  assign mem_MPORT_241_addr = 9'hf1;
  assign mem_MPORT_241_mask = 1'h1;
  assign mem_MPORT_241_en = reset;
  assign mem_MPORT_242_data = 19'h0;
  assign mem_MPORT_242_addr = 9'hf2;
  assign mem_MPORT_242_mask = 1'h1;
  assign mem_MPORT_242_en = reset;
  assign mem_MPORT_243_data = 19'h0;
  assign mem_MPORT_243_addr = 9'hf3;
  assign mem_MPORT_243_mask = 1'h1;
  assign mem_MPORT_243_en = reset;
  assign mem_MPORT_244_data = 19'h0;
  assign mem_MPORT_244_addr = 9'hf4;
  assign mem_MPORT_244_mask = 1'h1;
  assign mem_MPORT_244_en = reset;
  assign mem_MPORT_245_data = 19'h0;
  assign mem_MPORT_245_addr = 9'hf5;
  assign mem_MPORT_245_mask = 1'h1;
  assign mem_MPORT_245_en = reset;
  assign mem_MPORT_246_data = 19'h0;
  assign mem_MPORT_246_addr = 9'hf6;
  assign mem_MPORT_246_mask = 1'h1;
  assign mem_MPORT_246_en = reset;
  assign mem_MPORT_247_data = 19'h0;
  assign mem_MPORT_247_addr = 9'hf7;
  assign mem_MPORT_247_mask = 1'h1;
  assign mem_MPORT_247_en = reset;
  assign mem_MPORT_248_data = 19'h0;
  assign mem_MPORT_248_addr = 9'hf8;
  assign mem_MPORT_248_mask = 1'h1;
  assign mem_MPORT_248_en = reset;
  assign mem_MPORT_249_data = 19'h0;
  assign mem_MPORT_249_addr = 9'hf9;
  assign mem_MPORT_249_mask = 1'h1;
  assign mem_MPORT_249_en = reset;
  assign mem_MPORT_250_data = 19'h0;
  assign mem_MPORT_250_addr = 9'hfa;
  assign mem_MPORT_250_mask = 1'h1;
  assign mem_MPORT_250_en = reset;
  assign mem_MPORT_251_data = 19'h0;
  assign mem_MPORT_251_addr = 9'hfb;
  assign mem_MPORT_251_mask = 1'h1;
  assign mem_MPORT_251_en = reset;
  assign mem_MPORT_252_data = 19'h0;
  assign mem_MPORT_252_addr = 9'hfc;
  assign mem_MPORT_252_mask = 1'h1;
  assign mem_MPORT_252_en = reset;
  assign mem_MPORT_253_data = 19'h0;
  assign mem_MPORT_253_addr = 9'hfd;
  assign mem_MPORT_253_mask = 1'h1;
  assign mem_MPORT_253_en = reset;
  assign mem_MPORT_254_data = 19'h0;
  assign mem_MPORT_254_addr = 9'hfe;
  assign mem_MPORT_254_mask = 1'h1;
  assign mem_MPORT_254_en = reset;
  assign mem_MPORT_255_data = 19'h0;
  assign mem_MPORT_255_addr = 9'hff;
  assign mem_MPORT_255_mask = 1'h1;
  assign mem_MPORT_255_en = reset;
  assign mem_MPORT_256_data = 19'h0;
  assign mem_MPORT_256_addr = 9'h100;
  assign mem_MPORT_256_mask = 1'h1;
  assign mem_MPORT_256_en = reset;
  assign mem_MPORT_257_data = 19'h0;
  assign mem_MPORT_257_addr = 9'h101;
  assign mem_MPORT_257_mask = 1'h1;
  assign mem_MPORT_257_en = reset;
  assign mem_MPORT_258_data = 19'h0;
  assign mem_MPORT_258_addr = 9'h102;
  assign mem_MPORT_258_mask = 1'h1;
  assign mem_MPORT_258_en = reset;
  assign mem_MPORT_259_data = 19'h0;
  assign mem_MPORT_259_addr = 9'h103;
  assign mem_MPORT_259_mask = 1'h1;
  assign mem_MPORT_259_en = reset;
  assign mem_MPORT_260_data = 19'h0;
  assign mem_MPORT_260_addr = 9'h104;
  assign mem_MPORT_260_mask = 1'h1;
  assign mem_MPORT_260_en = reset;
  assign mem_MPORT_261_data = 19'h0;
  assign mem_MPORT_261_addr = 9'h105;
  assign mem_MPORT_261_mask = 1'h1;
  assign mem_MPORT_261_en = reset;
  assign mem_MPORT_262_data = 19'h0;
  assign mem_MPORT_262_addr = 9'h106;
  assign mem_MPORT_262_mask = 1'h1;
  assign mem_MPORT_262_en = reset;
  assign mem_MPORT_263_data = 19'h0;
  assign mem_MPORT_263_addr = 9'h107;
  assign mem_MPORT_263_mask = 1'h1;
  assign mem_MPORT_263_en = reset;
  assign mem_MPORT_264_data = 19'h0;
  assign mem_MPORT_264_addr = 9'h108;
  assign mem_MPORT_264_mask = 1'h1;
  assign mem_MPORT_264_en = reset;
  assign mem_MPORT_265_data = 19'h0;
  assign mem_MPORT_265_addr = 9'h109;
  assign mem_MPORT_265_mask = 1'h1;
  assign mem_MPORT_265_en = reset;
  assign mem_MPORT_266_data = 19'h0;
  assign mem_MPORT_266_addr = 9'h10a;
  assign mem_MPORT_266_mask = 1'h1;
  assign mem_MPORT_266_en = reset;
  assign mem_MPORT_267_data = 19'h0;
  assign mem_MPORT_267_addr = 9'h10b;
  assign mem_MPORT_267_mask = 1'h1;
  assign mem_MPORT_267_en = reset;
  assign mem_MPORT_268_data = 19'h0;
  assign mem_MPORT_268_addr = 9'h10c;
  assign mem_MPORT_268_mask = 1'h1;
  assign mem_MPORT_268_en = reset;
  assign mem_MPORT_269_data = 19'h0;
  assign mem_MPORT_269_addr = 9'h10d;
  assign mem_MPORT_269_mask = 1'h1;
  assign mem_MPORT_269_en = reset;
  assign mem_MPORT_270_data = 19'h0;
  assign mem_MPORT_270_addr = 9'h10e;
  assign mem_MPORT_270_mask = 1'h1;
  assign mem_MPORT_270_en = reset;
  assign mem_MPORT_271_data = 19'h0;
  assign mem_MPORT_271_addr = 9'h10f;
  assign mem_MPORT_271_mask = 1'h1;
  assign mem_MPORT_271_en = reset;
  assign mem_MPORT_272_data = 19'h0;
  assign mem_MPORT_272_addr = 9'h110;
  assign mem_MPORT_272_mask = 1'h1;
  assign mem_MPORT_272_en = reset;
  assign mem_MPORT_273_data = 19'h0;
  assign mem_MPORT_273_addr = 9'h111;
  assign mem_MPORT_273_mask = 1'h1;
  assign mem_MPORT_273_en = reset;
  assign mem_MPORT_274_data = 19'h0;
  assign mem_MPORT_274_addr = 9'h112;
  assign mem_MPORT_274_mask = 1'h1;
  assign mem_MPORT_274_en = reset;
  assign mem_MPORT_275_data = 19'h0;
  assign mem_MPORT_275_addr = 9'h113;
  assign mem_MPORT_275_mask = 1'h1;
  assign mem_MPORT_275_en = reset;
  assign mem_MPORT_276_data = 19'h0;
  assign mem_MPORT_276_addr = 9'h114;
  assign mem_MPORT_276_mask = 1'h1;
  assign mem_MPORT_276_en = reset;
  assign mem_MPORT_277_data = 19'h0;
  assign mem_MPORT_277_addr = 9'h115;
  assign mem_MPORT_277_mask = 1'h1;
  assign mem_MPORT_277_en = reset;
  assign mem_MPORT_278_data = 19'h0;
  assign mem_MPORT_278_addr = 9'h116;
  assign mem_MPORT_278_mask = 1'h1;
  assign mem_MPORT_278_en = reset;
  assign mem_MPORT_279_data = 19'h0;
  assign mem_MPORT_279_addr = 9'h117;
  assign mem_MPORT_279_mask = 1'h1;
  assign mem_MPORT_279_en = reset;
  assign mem_MPORT_280_data = 19'h0;
  assign mem_MPORT_280_addr = 9'h118;
  assign mem_MPORT_280_mask = 1'h1;
  assign mem_MPORT_280_en = reset;
  assign mem_MPORT_281_data = 19'h0;
  assign mem_MPORT_281_addr = 9'h119;
  assign mem_MPORT_281_mask = 1'h1;
  assign mem_MPORT_281_en = reset;
  assign mem_MPORT_282_data = 19'h0;
  assign mem_MPORT_282_addr = 9'h11a;
  assign mem_MPORT_282_mask = 1'h1;
  assign mem_MPORT_282_en = reset;
  assign mem_MPORT_283_data = 19'h0;
  assign mem_MPORT_283_addr = 9'h11b;
  assign mem_MPORT_283_mask = 1'h1;
  assign mem_MPORT_283_en = reset;
  assign mem_MPORT_284_data = 19'h0;
  assign mem_MPORT_284_addr = 9'h11c;
  assign mem_MPORT_284_mask = 1'h1;
  assign mem_MPORT_284_en = reset;
  assign mem_MPORT_285_data = 19'h0;
  assign mem_MPORT_285_addr = 9'h11d;
  assign mem_MPORT_285_mask = 1'h1;
  assign mem_MPORT_285_en = reset;
  assign mem_MPORT_286_data = 19'h0;
  assign mem_MPORT_286_addr = 9'h11e;
  assign mem_MPORT_286_mask = 1'h1;
  assign mem_MPORT_286_en = reset;
  assign mem_MPORT_287_data = 19'h0;
  assign mem_MPORT_287_addr = 9'h11f;
  assign mem_MPORT_287_mask = 1'h1;
  assign mem_MPORT_287_en = reset;
  assign mem_MPORT_288_data = 19'h0;
  assign mem_MPORT_288_addr = 9'h120;
  assign mem_MPORT_288_mask = 1'h1;
  assign mem_MPORT_288_en = reset;
  assign mem_MPORT_289_data = 19'h0;
  assign mem_MPORT_289_addr = 9'h121;
  assign mem_MPORT_289_mask = 1'h1;
  assign mem_MPORT_289_en = reset;
  assign mem_MPORT_290_data = 19'h0;
  assign mem_MPORT_290_addr = 9'h122;
  assign mem_MPORT_290_mask = 1'h1;
  assign mem_MPORT_290_en = reset;
  assign mem_MPORT_291_data = 19'h0;
  assign mem_MPORT_291_addr = 9'h123;
  assign mem_MPORT_291_mask = 1'h1;
  assign mem_MPORT_291_en = reset;
  assign mem_MPORT_292_data = 19'h0;
  assign mem_MPORT_292_addr = 9'h124;
  assign mem_MPORT_292_mask = 1'h1;
  assign mem_MPORT_292_en = reset;
  assign mem_MPORT_293_data = 19'h0;
  assign mem_MPORT_293_addr = 9'h125;
  assign mem_MPORT_293_mask = 1'h1;
  assign mem_MPORT_293_en = reset;
  assign mem_MPORT_294_data = 19'h0;
  assign mem_MPORT_294_addr = 9'h126;
  assign mem_MPORT_294_mask = 1'h1;
  assign mem_MPORT_294_en = reset;
  assign mem_MPORT_295_data = 19'h0;
  assign mem_MPORT_295_addr = 9'h127;
  assign mem_MPORT_295_mask = 1'h1;
  assign mem_MPORT_295_en = reset;
  assign mem_MPORT_296_data = 19'h0;
  assign mem_MPORT_296_addr = 9'h128;
  assign mem_MPORT_296_mask = 1'h1;
  assign mem_MPORT_296_en = reset;
  assign mem_MPORT_297_data = 19'h0;
  assign mem_MPORT_297_addr = 9'h129;
  assign mem_MPORT_297_mask = 1'h1;
  assign mem_MPORT_297_en = reset;
  assign mem_MPORT_298_data = 19'h0;
  assign mem_MPORT_298_addr = 9'h12a;
  assign mem_MPORT_298_mask = 1'h1;
  assign mem_MPORT_298_en = reset;
  assign mem_MPORT_299_data = 19'h0;
  assign mem_MPORT_299_addr = 9'h12b;
  assign mem_MPORT_299_mask = 1'h1;
  assign mem_MPORT_299_en = reset;
  assign mem_MPORT_300_data = 19'h0;
  assign mem_MPORT_300_addr = 9'h12c;
  assign mem_MPORT_300_mask = 1'h1;
  assign mem_MPORT_300_en = reset;
  assign mem_MPORT_301_data = 19'h0;
  assign mem_MPORT_301_addr = 9'h12d;
  assign mem_MPORT_301_mask = 1'h1;
  assign mem_MPORT_301_en = reset;
  assign mem_MPORT_302_data = 19'h0;
  assign mem_MPORT_302_addr = 9'h12e;
  assign mem_MPORT_302_mask = 1'h1;
  assign mem_MPORT_302_en = reset;
  assign mem_MPORT_303_data = 19'h0;
  assign mem_MPORT_303_addr = 9'h12f;
  assign mem_MPORT_303_mask = 1'h1;
  assign mem_MPORT_303_en = reset;
  assign mem_MPORT_304_data = 19'h0;
  assign mem_MPORT_304_addr = 9'h130;
  assign mem_MPORT_304_mask = 1'h1;
  assign mem_MPORT_304_en = reset;
  assign mem_MPORT_305_data = 19'h0;
  assign mem_MPORT_305_addr = 9'h131;
  assign mem_MPORT_305_mask = 1'h1;
  assign mem_MPORT_305_en = reset;
  assign mem_MPORT_306_data = 19'h0;
  assign mem_MPORT_306_addr = 9'h132;
  assign mem_MPORT_306_mask = 1'h1;
  assign mem_MPORT_306_en = reset;
  assign mem_MPORT_307_data = 19'h0;
  assign mem_MPORT_307_addr = 9'h133;
  assign mem_MPORT_307_mask = 1'h1;
  assign mem_MPORT_307_en = reset;
  assign mem_MPORT_308_data = 19'h0;
  assign mem_MPORT_308_addr = 9'h134;
  assign mem_MPORT_308_mask = 1'h1;
  assign mem_MPORT_308_en = reset;
  assign mem_MPORT_309_data = 19'h0;
  assign mem_MPORT_309_addr = 9'h135;
  assign mem_MPORT_309_mask = 1'h1;
  assign mem_MPORT_309_en = reset;
  assign mem_MPORT_310_data = 19'h0;
  assign mem_MPORT_310_addr = 9'h136;
  assign mem_MPORT_310_mask = 1'h1;
  assign mem_MPORT_310_en = reset;
  assign mem_MPORT_311_data = 19'h0;
  assign mem_MPORT_311_addr = 9'h137;
  assign mem_MPORT_311_mask = 1'h1;
  assign mem_MPORT_311_en = reset;
  assign mem_MPORT_312_data = 19'h0;
  assign mem_MPORT_312_addr = 9'h138;
  assign mem_MPORT_312_mask = 1'h1;
  assign mem_MPORT_312_en = reset;
  assign mem_MPORT_313_data = 19'h0;
  assign mem_MPORT_313_addr = 9'h139;
  assign mem_MPORT_313_mask = 1'h1;
  assign mem_MPORT_313_en = reset;
  assign mem_MPORT_314_data = 19'h0;
  assign mem_MPORT_314_addr = 9'h13a;
  assign mem_MPORT_314_mask = 1'h1;
  assign mem_MPORT_314_en = reset;
  assign mem_MPORT_315_data = 19'h0;
  assign mem_MPORT_315_addr = 9'h13b;
  assign mem_MPORT_315_mask = 1'h1;
  assign mem_MPORT_315_en = reset;
  assign mem_MPORT_316_data = 19'h0;
  assign mem_MPORT_316_addr = 9'h13c;
  assign mem_MPORT_316_mask = 1'h1;
  assign mem_MPORT_316_en = reset;
  assign mem_MPORT_317_data = 19'h0;
  assign mem_MPORT_317_addr = 9'h13d;
  assign mem_MPORT_317_mask = 1'h1;
  assign mem_MPORT_317_en = reset;
  assign mem_MPORT_318_data = 19'h0;
  assign mem_MPORT_318_addr = 9'h13e;
  assign mem_MPORT_318_mask = 1'h1;
  assign mem_MPORT_318_en = reset;
  assign mem_MPORT_319_data = 19'h0;
  assign mem_MPORT_319_addr = 9'h13f;
  assign mem_MPORT_319_mask = 1'h1;
  assign mem_MPORT_319_en = reset;
  assign mem_MPORT_320_data = 19'h0;
  assign mem_MPORT_320_addr = 9'h140;
  assign mem_MPORT_320_mask = 1'h1;
  assign mem_MPORT_320_en = reset;
  assign mem_MPORT_321_data = 19'h0;
  assign mem_MPORT_321_addr = 9'h141;
  assign mem_MPORT_321_mask = 1'h1;
  assign mem_MPORT_321_en = reset;
  assign mem_MPORT_322_data = 19'h0;
  assign mem_MPORT_322_addr = 9'h142;
  assign mem_MPORT_322_mask = 1'h1;
  assign mem_MPORT_322_en = reset;
  assign mem_MPORT_323_data = 19'h0;
  assign mem_MPORT_323_addr = 9'h143;
  assign mem_MPORT_323_mask = 1'h1;
  assign mem_MPORT_323_en = reset;
  assign mem_MPORT_324_data = 19'h0;
  assign mem_MPORT_324_addr = 9'h144;
  assign mem_MPORT_324_mask = 1'h1;
  assign mem_MPORT_324_en = reset;
  assign mem_MPORT_325_data = 19'h0;
  assign mem_MPORT_325_addr = 9'h145;
  assign mem_MPORT_325_mask = 1'h1;
  assign mem_MPORT_325_en = reset;
  assign mem_MPORT_326_data = 19'h0;
  assign mem_MPORT_326_addr = 9'h146;
  assign mem_MPORT_326_mask = 1'h1;
  assign mem_MPORT_326_en = reset;
  assign mem_MPORT_327_data = 19'h0;
  assign mem_MPORT_327_addr = 9'h147;
  assign mem_MPORT_327_mask = 1'h1;
  assign mem_MPORT_327_en = reset;
  assign mem_MPORT_328_data = 19'h0;
  assign mem_MPORT_328_addr = 9'h148;
  assign mem_MPORT_328_mask = 1'h1;
  assign mem_MPORT_328_en = reset;
  assign mem_MPORT_329_data = 19'h0;
  assign mem_MPORT_329_addr = 9'h149;
  assign mem_MPORT_329_mask = 1'h1;
  assign mem_MPORT_329_en = reset;
  assign mem_MPORT_330_data = 19'h0;
  assign mem_MPORT_330_addr = 9'h14a;
  assign mem_MPORT_330_mask = 1'h1;
  assign mem_MPORT_330_en = reset;
  assign mem_MPORT_331_data = 19'h0;
  assign mem_MPORT_331_addr = 9'h14b;
  assign mem_MPORT_331_mask = 1'h1;
  assign mem_MPORT_331_en = reset;
  assign mem_MPORT_332_data = 19'h0;
  assign mem_MPORT_332_addr = 9'h14c;
  assign mem_MPORT_332_mask = 1'h1;
  assign mem_MPORT_332_en = reset;
  assign mem_MPORT_333_data = 19'h0;
  assign mem_MPORT_333_addr = 9'h14d;
  assign mem_MPORT_333_mask = 1'h1;
  assign mem_MPORT_333_en = reset;
  assign mem_MPORT_334_data = 19'h0;
  assign mem_MPORT_334_addr = 9'h14e;
  assign mem_MPORT_334_mask = 1'h1;
  assign mem_MPORT_334_en = reset;
  assign mem_MPORT_335_data = 19'h0;
  assign mem_MPORT_335_addr = 9'h14f;
  assign mem_MPORT_335_mask = 1'h1;
  assign mem_MPORT_335_en = reset;
  assign mem_MPORT_336_data = 19'h0;
  assign mem_MPORT_336_addr = 9'h150;
  assign mem_MPORT_336_mask = 1'h1;
  assign mem_MPORT_336_en = reset;
  assign mem_MPORT_337_data = 19'h0;
  assign mem_MPORT_337_addr = 9'h151;
  assign mem_MPORT_337_mask = 1'h1;
  assign mem_MPORT_337_en = reset;
  assign mem_MPORT_338_data = 19'h0;
  assign mem_MPORT_338_addr = 9'h152;
  assign mem_MPORT_338_mask = 1'h1;
  assign mem_MPORT_338_en = reset;
  assign mem_MPORT_339_data = 19'h0;
  assign mem_MPORT_339_addr = 9'h153;
  assign mem_MPORT_339_mask = 1'h1;
  assign mem_MPORT_339_en = reset;
  assign mem_MPORT_340_data = 19'h0;
  assign mem_MPORT_340_addr = 9'h154;
  assign mem_MPORT_340_mask = 1'h1;
  assign mem_MPORT_340_en = reset;
  assign mem_MPORT_341_data = 19'h0;
  assign mem_MPORT_341_addr = 9'h155;
  assign mem_MPORT_341_mask = 1'h1;
  assign mem_MPORT_341_en = reset;
  assign mem_MPORT_342_data = 19'h0;
  assign mem_MPORT_342_addr = 9'h156;
  assign mem_MPORT_342_mask = 1'h1;
  assign mem_MPORT_342_en = reset;
  assign mem_MPORT_343_data = 19'h0;
  assign mem_MPORT_343_addr = 9'h157;
  assign mem_MPORT_343_mask = 1'h1;
  assign mem_MPORT_343_en = reset;
  assign mem_MPORT_344_data = 19'h0;
  assign mem_MPORT_344_addr = 9'h158;
  assign mem_MPORT_344_mask = 1'h1;
  assign mem_MPORT_344_en = reset;
  assign mem_MPORT_345_data = 19'h0;
  assign mem_MPORT_345_addr = 9'h159;
  assign mem_MPORT_345_mask = 1'h1;
  assign mem_MPORT_345_en = reset;
  assign mem_MPORT_346_data = 19'h0;
  assign mem_MPORT_346_addr = 9'h15a;
  assign mem_MPORT_346_mask = 1'h1;
  assign mem_MPORT_346_en = reset;
  assign mem_MPORT_347_data = 19'h0;
  assign mem_MPORT_347_addr = 9'h15b;
  assign mem_MPORT_347_mask = 1'h1;
  assign mem_MPORT_347_en = reset;
  assign mem_MPORT_348_data = 19'h0;
  assign mem_MPORT_348_addr = 9'h15c;
  assign mem_MPORT_348_mask = 1'h1;
  assign mem_MPORT_348_en = reset;
  assign mem_MPORT_349_data = 19'h0;
  assign mem_MPORT_349_addr = 9'h15d;
  assign mem_MPORT_349_mask = 1'h1;
  assign mem_MPORT_349_en = reset;
  assign mem_MPORT_350_data = 19'h0;
  assign mem_MPORT_350_addr = 9'h15e;
  assign mem_MPORT_350_mask = 1'h1;
  assign mem_MPORT_350_en = reset;
  assign mem_MPORT_351_data = 19'h0;
  assign mem_MPORT_351_addr = 9'h15f;
  assign mem_MPORT_351_mask = 1'h1;
  assign mem_MPORT_351_en = reset;
  assign mem_MPORT_352_data = 19'h0;
  assign mem_MPORT_352_addr = 9'h160;
  assign mem_MPORT_352_mask = 1'h1;
  assign mem_MPORT_352_en = reset;
  assign mem_MPORT_353_data = 19'h0;
  assign mem_MPORT_353_addr = 9'h161;
  assign mem_MPORT_353_mask = 1'h1;
  assign mem_MPORT_353_en = reset;
  assign mem_MPORT_354_data = 19'h0;
  assign mem_MPORT_354_addr = 9'h162;
  assign mem_MPORT_354_mask = 1'h1;
  assign mem_MPORT_354_en = reset;
  assign mem_MPORT_355_data = 19'h0;
  assign mem_MPORT_355_addr = 9'h163;
  assign mem_MPORT_355_mask = 1'h1;
  assign mem_MPORT_355_en = reset;
  assign mem_MPORT_356_data = 19'h0;
  assign mem_MPORT_356_addr = 9'h164;
  assign mem_MPORT_356_mask = 1'h1;
  assign mem_MPORT_356_en = reset;
  assign mem_MPORT_357_data = 19'h0;
  assign mem_MPORT_357_addr = 9'h165;
  assign mem_MPORT_357_mask = 1'h1;
  assign mem_MPORT_357_en = reset;
  assign mem_MPORT_358_data = 19'h0;
  assign mem_MPORT_358_addr = 9'h166;
  assign mem_MPORT_358_mask = 1'h1;
  assign mem_MPORT_358_en = reset;
  assign mem_MPORT_359_data = 19'h0;
  assign mem_MPORT_359_addr = 9'h167;
  assign mem_MPORT_359_mask = 1'h1;
  assign mem_MPORT_359_en = reset;
  assign mem_MPORT_360_data = 19'h0;
  assign mem_MPORT_360_addr = 9'h168;
  assign mem_MPORT_360_mask = 1'h1;
  assign mem_MPORT_360_en = reset;
  assign mem_MPORT_361_data = 19'h0;
  assign mem_MPORT_361_addr = 9'h169;
  assign mem_MPORT_361_mask = 1'h1;
  assign mem_MPORT_361_en = reset;
  assign mem_MPORT_362_data = 19'h0;
  assign mem_MPORT_362_addr = 9'h16a;
  assign mem_MPORT_362_mask = 1'h1;
  assign mem_MPORT_362_en = reset;
  assign mem_MPORT_363_data = 19'h0;
  assign mem_MPORT_363_addr = 9'h16b;
  assign mem_MPORT_363_mask = 1'h1;
  assign mem_MPORT_363_en = reset;
  assign mem_MPORT_364_data = 19'h0;
  assign mem_MPORT_364_addr = 9'h16c;
  assign mem_MPORT_364_mask = 1'h1;
  assign mem_MPORT_364_en = reset;
  assign mem_MPORT_365_data = 19'h0;
  assign mem_MPORT_365_addr = 9'h16d;
  assign mem_MPORT_365_mask = 1'h1;
  assign mem_MPORT_365_en = reset;
  assign mem_MPORT_366_data = 19'h0;
  assign mem_MPORT_366_addr = 9'h16e;
  assign mem_MPORT_366_mask = 1'h1;
  assign mem_MPORT_366_en = reset;
  assign mem_MPORT_367_data = 19'h0;
  assign mem_MPORT_367_addr = 9'h16f;
  assign mem_MPORT_367_mask = 1'h1;
  assign mem_MPORT_367_en = reset;
  assign mem_MPORT_368_data = 19'h0;
  assign mem_MPORT_368_addr = 9'h170;
  assign mem_MPORT_368_mask = 1'h1;
  assign mem_MPORT_368_en = reset;
  assign mem_MPORT_369_data = 19'h0;
  assign mem_MPORT_369_addr = 9'h171;
  assign mem_MPORT_369_mask = 1'h1;
  assign mem_MPORT_369_en = reset;
  assign mem_MPORT_370_data = 19'h0;
  assign mem_MPORT_370_addr = 9'h172;
  assign mem_MPORT_370_mask = 1'h1;
  assign mem_MPORT_370_en = reset;
  assign mem_MPORT_371_data = 19'h0;
  assign mem_MPORT_371_addr = 9'h173;
  assign mem_MPORT_371_mask = 1'h1;
  assign mem_MPORT_371_en = reset;
  assign mem_MPORT_372_data = 19'h0;
  assign mem_MPORT_372_addr = 9'h174;
  assign mem_MPORT_372_mask = 1'h1;
  assign mem_MPORT_372_en = reset;
  assign mem_MPORT_373_data = 19'h0;
  assign mem_MPORT_373_addr = 9'h175;
  assign mem_MPORT_373_mask = 1'h1;
  assign mem_MPORT_373_en = reset;
  assign mem_MPORT_374_data = 19'h0;
  assign mem_MPORT_374_addr = 9'h176;
  assign mem_MPORT_374_mask = 1'h1;
  assign mem_MPORT_374_en = reset;
  assign mem_MPORT_375_data = 19'h0;
  assign mem_MPORT_375_addr = 9'h177;
  assign mem_MPORT_375_mask = 1'h1;
  assign mem_MPORT_375_en = reset;
  assign mem_MPORT_376_data = 19'h0;
  assign mem_MPORT_376_addr = 9'h178;
  assign mem_MPORT_376_mask = 1'h1;
  assign mem_MPORT_376_en = reset;
  assign mem_MPORT_377_data = 19'h0;
  assign mem_MPORT_377_addr = 9'h179;
  assign mem_MPORT_377_mask = 1'h1;
  assign mem_MPORT_377_en = reset;
  assign mem_MPORT_378_data = 19'h0;
  assign mem_MPORT_378_addr = 9'h17a;
  assign mem_MPORT_378_mask = 1'h1;
  assign mem_MPORT_378_en = reset;
  assign mem_MPORT_379_data = 19'h0;
  assign mem_MPORT_379_addr = 9'h17b;
  assign mem_MPORT_379_mask = 1'h1;
  assign mem_MPORT_379_en = reset;
  assign mem_MPORT_380_data = 19'h0;
  assign mem_MPORT_380_addr = 9'h17c;
  assign mem_MPORT_380_mask = 1'h1;
  assign mem_MPORT_380_en = reset;
  assign mem_MPORT_381_data = 19'h0;
  assign mem_MPORT_381_addr = 9'h17d;
  assign mem_MPORT_381_mask = 1'h1;
  assign mem_MPORT_381_en = reset;
  assign mem_MPORT_382_data = 19'h0;
  assign mem_MPORT_382_addr = 9'h17e;
  assign mem_MPORT_382_mask = 1'h1;
  assign mem_MPORT_382_en = reset;
  assign mem_MPORT_383_data = 19'h0;
  assign mem_MPORT_383_addr = 9'h17f;
  assign mem_MPORT_383_mask = 1'h1;
  assign mem_MPORT_383_en = reset;
  assign mem_MPORT_384_data = 19'h0;
  assign mem_MPORT_384_addr = 9'h180;
  assign mem_MPORT_384_mask = 1'h1;
  assign mem_MPORT_384_en = reset;
  assign mem_MPORT_385_data = 19'h0;
  assign mem_MPORT_385_addr = 9'h181;
  assign mem_MPORT_385_mask = 1'h1;
  assign mem_MPORT_385_en = reset;
  assign mem_MPORT_386_data = 19'h0;
  assign mem_MPORT_386_addr = 9'h182;
  assign mem_MPORT_386_mask = 1'h1;
  assign mem_MPORT_386_en = reset;
  assign mem_MPORT_387_data = 19'h0;
  assign mem_MPORT_387_addr = 9'h183;
  assign mem_MPORT_387_mask = 1'h1;
  assign mem_MPORT_387_en = reset;
  assign mem_MPORT_388_data = 19'h0;
  assign mem_MPORT_388_addr = 9'h184;
  assign mem_MPORT_388_mask = 1'h1;
  assign mem_MPORT_388_en = reset;
  assign mem_MPORT_389_data = 19'h0;
  assign mem_MPORT_389_addr = 9'h185;
  assign mem_MPORT_389_mask = 1'h1;
  assign mem_MPORT_389_en = reset;
  assign mem_MPORT_390_data = 19'h0;
  assign mem_MPORT_390_addr = 9'h186;
  assign mem_MPORT_390_mask = 1'h1;
  assign mem_MPORT_390_en = reset;
  assign mem_MPORT_391_data = 19'h0;
  assign mem_MPORT_391_addr = 9'h187;
  assign mem_MPORT_391_mask = 1'h1;
  assign mem_MPORT_391_en = reset;
  assign mem_MPORT_392_data = 19'h0;
  assign mem_MPORT_392_addr = 9'h188;
  assign mem_MPORT_392_mask = 1'h1;
  assign mem_MPORT_392_en = reset;
  assign mem_MPORT_393_data = 19'h0;
  assign mem_MPORT_393_addr = 9'h189;
  assign mem_MPORT_393_mask = 1'h1;
  assign mem_MPORT_393_en = reset;
  assign mem_MPORT_394_data = 19'h0;
  assign mem_MPORT_394_addr = 9'h18a;
  assign mem_MPORT_394_mask = 1'h1;
  assign mem_MPORT_394_en = reset;
  assign mem_MPORT_395_data = 19'h0;
  assign mem_MPORT_395_addr = 9'h18b;
  assign mem_MPORT_395_mask = 1'h1;
  assign mem_MPORT_395_en = reset;
  assign mem_MPORT_396_data = 19'h0;
  assign mem_MPORT_396_addr = 9'h18c;
  assign mem_MPORT_396_mask = 1'h1;
  assign mem_MPORT_396_en = reset;
  assign mem_MPORT_397_data = 19'h0;
  assign mem_MPORT_397_addr = 9'h18d;
  assign mem_MPORT_397_mask = 1'h1;
  assign mem_MPORT_397_en = reset;
  assign mem_MPORT_398_data = 19'h0;
  assign mem_MPORT_398_addr = 9'h18e;
  assign mem_MPORT_398_mask = 1'h1;
  assign mem_MPORT_398_en = reset;
  assign mem_MPORT_399_data = 19'h0;
  assign mem_MPORT_399_addr = 9'h18f;
  assign mem_MPORT_399_mask = 1'h1;
  assign mem_MPORT_399_en = reset;
  assign mem_MPORT_400_data = 19'h0;
  assign mem_MPORT_400_addr = 9'h190;
  assign mem_MPORT_400_mask = 1'h1;
  assign mem_MPORT_400_en = reset;
  assign mem_MPORT_401_data = 19'h0;
  assign mem_MPORT_401_addr = 9'h191;
  assign mem_MPORT_401_mask = 1'h1;
  assign mem_MPORT_401_en = reset;
  assign mem_MPORT_402_data = 19'h0;
  assign mem_MPORT_402_addr = 9'h192;
  assign mem_MPORT_402_mask = 1'h1;
  assign mem_MPORT_402_en = reset;
  assign mem_MPORT_403_data = 19'h0;
  assign mem_MPORT_403_addr = 9'h193;
  assign mem_MPORT_403_mask = 1'h1;
  assign mem_MPORT_403_en = reset;
  assign mem_MPORT_404_data = 19'h0;
  assign mem_MPORT_404_addr = 9'h194;
  assign mem_MPORT_404_mask = 1'h1;
  assign mem_MPORT_404_en = reset;
  assign mem_MPORT_405_data = 19'h0;
  assign mem_MPORT_405_addr = 9'h195;
  assign mem_MPORT_405_mask = 1'h1;
  assign mem_MPORT_405_en = reset;
  assign mem_MPORT_406_data = 19'h0;
  assign mem_MPORT_406_addr = 9'h196;
  assign mem_MPORT_406_mask = 1'h1;
  assign mem_MPORT_406_en = reset;
  assign mem_MPORT_407_data = 19'h0;
  assign mem_MPORT_407_addr = 9'h197;
  assign mem_MPORT_407_mask = 1'h1;
  assign mem_MPORT_407_en = reset;
  assign mem_MPORT_408_data = 19'h0;
  assign mem_MPORT_408_addr = 9'h198;
  assign mem_MPORT_408_mask = 1'h1;
  assign mem_MPORT_408_en = reset;
  assign mem_MPORT_409_data = 19'h0;
  assign mem_MPORT_409_addr = 9'h199;
  assign mem_MPORT_409_mask = 1'h1;
  assign mem_MPORT_409_en = reset;
  assign mem_MPORT_410_data = 19'h0;
  assign mem_MPORT_410_addr = 9'h19a;
  assign mem_MPORT_410_mask = 1'h1;
  assign mem_MPORT_410_en = reset;
  assign mem_MPORT_411_data = 19'h0;
  assign mem_MPORT_411_addr = 9'h19b;
  assign mem_MPORT_411_mask = 1'h1;
  assign mem_MPORT_411_en = reset;
  assign mem_MPORT_412_data = 19'h0;
  assign mem_MPORT_412_addr = 9'h19c;
  assign mem_MPORT_412_mask = 1'h1;
  assign mem_MPORT_412_en = reset;
  assign mem_MPORT_413_data = 19'h0;
  assign mem_MPORT_413_addr = 9'h19d;
  assign mem_MPORT_413_mask = 1'h1;
  assign mem_MPORT_413_en = reset;
  assign mem_MPORT_414_data = 19'h0;
  assign mem_MPORT_414_addr = 9'h19e;
  assign mem_MPORT_414_mask = 1'h1;
  assign mem_MPORT_414_en = reset;
  assign mem_MPORT_415_data = 19'h0;
  assign mem_MPORT_415_addr = 9'h19f;
  assign mem_MPORT_415_mask = 1'h1;
  assign mem_MPORT_415_en = reset;
  assign mem_MPORT_416_data = 19'h0;
  assign mem_MPORT_416_addr = 9'h1a0;
  assign mem_MPORT_416_mask = 1'h1;
  assign mem_MPORT_416_en = reset;
  assign mem_MPORT_417_data = 19'h0;
  assign mem_MPORT_417_addr = 9'h1a1;
  assign mem_MPORT_417_mask = 1'h1;
  assign mem_MPORT_417_en = reset;
  assign mem_MPORT_418_data = 19'h0;
  assign mem_MPORT_418_addr = 9'h1a2;
  assign mem_MPORT_418_mask = 1'h1;
  assign mem_MPORT_418_en = reset;
  assign mem_MPORT_419_data = 19'h0;
  assign mem_MPORT_419_addr = 9'h1a3;
  assign mem_MPORT_419_mask = 1'h1;
  assign mem_MPORT_419_en = reset;
  assign mem_MPORT_420_data = 19'h0;
  assign mem_MPORT_420_addr = 9'h1a4;
  assign mem_MPORT_420_mask = 1'h1;
  assign mem_MPORT_420_en = reset;
  assign mem_MPORT_421_data = 19'h0;
  assign mem_MPORT_421_addr = 9'h1a5;
  assign mem_MPORT_421_mask = 1'h1;
  assign mem_MPORT_421_en = reset;
  assign mem_MPORT_422_data = 19'h0;
  assign mem_MPORT_422_addr = 9'h1a6;
  assign mem_MPORT_422_mask = 1'h1;
  assign mem_MPORT_422_en = reset;
  assign mem_MPORT_423_data = 19'h0;
  assign mem_MPORT_423_addr = 9'h1a7;
  assign mem_MPORT_423_mask = 1'h1;
  assign mem_MPORT_423_en = reset;
  assign mem_MPORT_424_data = 19'h0;
  assign mem_MPORT_424_addr = 9'h1a8;
  assign mem_MPORT_424_mask = 1'h1;
  assign mem_MPORT_424_en = reset;
  assign mem_MPORT_425_data = 19'h0;
  assign mem_MPORT_425_addr = 9'h1a9;
  assign mem_MPORT_425_mask = 1'h1;
  assign mem_MPORT_425_en = reset;
  assign mem_MPORT_426_data = 19'h0;
  assign mem_MPORT_426_addr = 9'h1aa;
  assign mem_MPORT_426_mask = 1'h1;
  assign mem_MPORT_426_en = reset;
  assign mem_MPORT_427_data = 19'h0;
  assign mem_MPORT_427_addr = 9'h1ab;
  assign mem_MPORT_427_mask = 1'h1;
  assign mem_MPORT_427_en = reset;
  assign mem_MPORT_428_data = 19'h0;
  assign mem_MPORT_428_addr = 9'h1ac;
  assign mem_MPORT_428_mask = 1'h1;
  assign mem_MPORT_428_en = reset;
  assign mem_MPORT_429_data = 19'h0;
  assign mem_MPORT_429_addr = 9'h1ad;
  assign mem_MPORT_429_mask = 1'h1;
  assign mem_MPORT_429_en = reset;
  assign mem_MPORT_430_data = 19'h0;
  assign mem_MPORT_430_addr = 9'h1ae;
  assign mem_MPORT_430_mask = 1'h1;
  assign mem_MPORT_430_en = reset;
  assign mem_MPORT_431_data = 19'h0;
  assign mem_MPORT_431_addr = 9'h1af;
  assign mem_MPORT_431_mask = 1'h1;
  assign mem_MPORT_431_en = reset;
  assign mem_MPORT_432_data = 19'h0;
  assign mem_MPORT_432_addr = 9'h1b0;
  assign mem_MPORT_432_mask = 1'h1;
  assign mem_MPORT_432_en = reset;
  assign mem_MPORT_433_data = 19'h0;
  assign mem_MPORT_433_addr = 9'h1b1;
  assign mem_MPORT_433_mask = 1'h1;
  assign mem_MPORT_433_en = reset;
  assign mem_MPORT_434_data = 19'h0;
  assign mem_MPORT_434_addr = 9'h1b2;
  assign mem_MPORT_434_mask = 1'h1;
  assign mem_MPORT_434_en = reset;
  assign mem_MPORT_435_data = 19'h0;
  assign mem_MPORT_435_addr = 9'h1b3;
  assign mem_MPORT_435_mask = 1'h1;
  assign mem_MPORT_435_en = reset;
  assign mem_MPORT_436_data = 19'h0;
  assign mem_MPORT_436_addr = 9'h1b4;
  assign mem_MPORT_436_mask = 1'h1;
  assign mem_MPORT_436_en = reset;
  assign mem_MPORT_437_data = 19'h0;
  assign mem_MPORT_437_addr = 9'h1b5;
  assign mem_MPORT_437_mask = 1'h1;
  assign mem_MPORT_437_en = reset;
  assign mem_MPORT_438_data = 19'h0;
  assign mem_MPORT_438_addr = 9'h1b6;
  assign mem_MPORT_438_mask = 1'h1;
  assign mem_MPORT_438_en = reset;
  assign mem_MPORT_439_data = 19'h0;
  assign mem_MPORT_439_addr = 9'h1b7;
  assign mem_MPORT_439_mask = 1'h1;
  assign mem_MPORT_439_en = reset;
  assign mem_MPORT_440_data = 19'h0;
  assign mem_MPORT_440_addr = 9'h1b8;
  assign mem_MPORT_440_mask = 1'h1;
  assign mem_MPORT_440_en = reset;
  assign mem_MPORT_441_data = 19'h0;
  assign mem_MPORT_441_addr = 9'h1b9;
  assign mem_MPORT_441_mask = 1'h1;
  assign mem_MPORT_441_en = reset;
  assign mem_MPORT_442_data = 19'h0;
  assign mem_MPORT_442_addr = 9'h1ba;
  assign mem_MPORT_442_mask = 1'h1;
  assign mem_MPORT_442_en = reset;
  assign mem_MPORT_443_data = 19'h0;
  assign mem_MPORT_443_addr = 9'h1bb;
  assign mem_MPORT_443_mask = 1'h1;
  assign mem_MPORT_443_en = reset;
  assign mem_MPORT_444_data = 19'h0;
  assign mem_MPORT_444_addr = 9'h1bc;
  assign mem_MPORT_444_mask = 1'h1;
  assign mem_MPORT_444_en = reset;
  assign mem_MPORT_445_data = 19'h0;
  assign mem_MPORT_445_addr = 9'h1bd;
  assign mem_MPORT_445_mask = 1'h1;
  assign mem_MPORT_445_en = reset;
  assign mem_MPORT_446_data = 19'h0;
  assign mem_MPORT_446_addr = 9'h1be;
  assign mem_MPORT_446_mask = 1'h1;
  assign mem_MPORT_446_en = reset;
  assign mem_MPORT_447_data = 19'h0;
  assign mem_MPORT_447_addr = 9'h1bf;
  assign mem_MPORT_447_mask = 1'h1;
  assign mem_MPORT_447_en = reset;
  assign mem_MPORT_448_data = 19'h0;
  assign mem_MPORT_448_addr = 9'h1c0;
  assign mem_MPORT_448_mask = 1'h1;
  assign mem_MPORT_448_en = reset;
  assign mem_MPORT_449_data = 19'h0;
  assign mem_MPORT_449_addr = 9'h1c1;
  assign mem_MPORT_449_mask = 1'h1;
  assign mem_MPORT_449_en = reset;
  assign mem_MPORT_450_data = 19'h0;
  assign mem_MPORT_450_addr = 9'h1c2;
  assign mem_MPORT_450_mask = 1'h1;
  assign mem_MPORT_450_en = reset;
  assign mem_MPORT_451_data = 19'h0;
  assign mem_MPORT_451_addr = 9'h1c3;
  assign mem_MPORT_451_mask = 1'h1;
  assign mem_MPORT_451_en = reset;
  assign mem_MPORT_452_data = 19'h0;
  assign mem_MPORT_452_addr = 9'h1c4;
  assign mem_MPORT_452_mask = 1'h1;
  assign mem_MPORT_452_en = reset;
  assign mem_MPORT_453_data = 19'h0;
  assign mem_MPORT_453_addr = 9'h1c5;
  assign mem_MPORT_453_mask = 1'h1;
  assign mem_MPORT_453_en = reset;
  assign mem_MPORT_454_data = 19'h0;
  assign mem_MPORT_454_addr = 9'h1c6;
  assign mem_MPORT_454_mask = 1'h1;
  assign mem_MPORT_454_en = reset;
  assign mem_MPORT_455_data = 19'h0;
  assign mem_MPORT_455_addr = 9'h1c7;
  assign mem_MPORT_455_mask = 1'h1;
  assign mem_MPORT_455_en = reset;
  assign mem_MPORT_456_data = 19'h0;
  assign mem_MPORT_456_addr = 9'h1c8;
  assign mem_MPORT_456_mask = 1'h1;
  assign mem_MPORT_456_en = reset;
  assign mem_MPORT_457_data = 19'h0;
  assign mem_MPORT_457_addr = 9'h1c9;
  assign mem_MPORT_457_mask = 1'h1;
  assign mem_MPORT_457_en = reset;
  assign mem_MPORT_458_data = 19'h0;
  assign mem_MPORT_458_addr = 9'h1ca;
  assign mem_MPORT_458_mask = 1'h1;
  assign mem_MPORT_458_en = reset;
  assign mem_MPORT_459_data = 19'h0;
  assign mem_MPORT_459_addr = 9'h1cb;
  assign mem_MPORT_459_mask = 1'h1;
  assign mem_MPORT_459_en = reset;
  assign mem_MPORT_460_data = 19'h0;
  assign mem_MPORT_460_addr = 9'h1cc;
  assign mem_MPORT_460_mask = 1'h1;
  assign mem_MPORT_460_en = reset;
  assign mem_MPORT_461_data = 19'h0;
  assign mem_MPORT_461_addr = 9'h1cd;
  assign mem_MPORT_461_mask = 1'h1;
  assign mem_MPORT_461_en = reset;
  assign mem_MPORT_462_data = 19'h0;
  assign mem_MPORT_462_addr = 9'h1ce;
  assign mem_MPORT_462_mask = 1'h1;
  assign mem_MPORT_462_en = reset;
  assign mem_MPORT_463_data = 19'h0;
  assign mem_MPORT_463_addr = 9'h1cf;
  assign mem_MPORT_463_mask = 1'h1;
  assign mem_MPORT_463_en = reset;
  assign mem_MPORT_464_data = 19'h0;
  assign mem_MPORT_464_addr = 9'h1d0;
  assign mem_MPORT_464_mask = 1'h1;
  assign mem_MPORT_464_en = reset;
  assign mem_MPORT_465_data = 19'h0;
  assign mem_MPORT_465_addr = 9'h1d1;
  assign mem_MPORT_465_mask = 1'h1;
  assign mem_MPORT_465_en = reset;
  assign mem_MPORT_466_data = 19'h0;
  assign mem_MPORT_466_addr = 9'h1d2;
  assign mem_MPORT_466_mask = 1'h1;
  assign mem_MPORT_466_en = reset;
  assign mem_MPORT_467_data = 19'h0;
  assign mem_MPORT_467_addr = 9'h1d3;
  assign mem_MPORT_467_mask = 1'h1;
  assign mem_MPORT_467_en = reset;
  assign mem_MPORT_468_data = 19'h0;
  assign mem_MPORT_468_addr = 9'h1d4;
  assign mem_MPORT_468_mask = 1'h1;
  assign mem_MPORT_468_en = reset;
  assign mem_MPORT_469_data = 19'h0;
  assign mem_MPORT_469_addr = 9'h1d5;
  assign mem_MPORT_469_mask = 1'h1;
  assign mem_MPORT_469_en = reset;
  assign mem_MPORT_470_data = 19'h0;
  assign mem_MPORT_470_addr = 9'h1d6;
  assign mem_MPORT_470_mask = 1'h1;
  assign mem_MPORT_470_en = reset;
  assign mem_MPORT_471_data = 19'h0;
  assign mem_MPORT_471_addr = 9'h1d7;
  assign mem_MPORT_471_mask = 1'h1;
  assign mem_MPORT_471_en = reset;
  assign mem_MPORT_472_data = 19'h0;
  assign mem_MPORT_472_addr = 9'h1d8;
  assign mem_MPORT_472_mask = 1'h1;
  assign mem_MPORT_472_en = reset;
  assign mem_MPORT_473_data = 19'h0;
  assign mem_MPORT_473_addr = 9'h1d9;
  assign mem_MPORT_473_mask = 1'h1;
  assign mem_MPORT_473_en = reset;
  assign mem_MPORT_474_data = 19'h0;
  assign mem_MPORT_474_addr = 9'h1da;
  assign mem_MPORT_474_mask = 1'h1;
  assign mem_MPORT_474_en = reset;
  assign mem_MPORT_475_data = 19'h0;
  assign mem_MPORT_475_addr = 9'h1db;
  assign mem_MPORT_475_mask = 1'h1;
  assign mem_MPORT_475_en = reset;
  assign mem_MPORT_476_data = 19'h0;
  assign mem_MPORT_476_addr = 9'h1dc;
  assign mem_MPORT_476_mask = 1'h1;
  assign mem_MPORT_476_en = reset;
  assign mem_MPORT_477_data = 19'h0;
  assign mem_MPORT_477_addr = 9'h1dd;
  assign mem_MPORT_477_mask = 1'h1;
  assign mem_MPORT_477_en = reset;
  assign mem_MPORT_478_data = 19'h0;
  assign mem_MPORT_478_addr = 9'h1de;
  assign mem_MPORT_478_mask = 1'h1;
  assign mem_MPORT_478_en = reset;
  assign mem_MPORT_479_data = 19'h0;
  assign mem_MPORT_479_addr = 9'h1df;
  assign mem_MPORT_479_mask = 1'h1;
  assign mem_MPORT_479_en = reset;
  assign mem_MPORT_480_data = 19'h0;
  assign mem_MPORT_480_addr = 9'h1e0;
  assign mem_MPORT_480_mask = 1'h1;
  assign mem_MPORT_480_en = reset;
  assign mem_MPORT_481_data = 19'h0;
  assign mem_MPORT_481_addr = 9'h1e1;
  assign mem_MPORT_481_mask = 1'h1;
  assign mem_MPORT_481_en = reset;
  assign mem_MPORT_482_data = 19'h0;
  assign mem_MPORT_482_addr = 9'h1e2;
  assign mem_MPORT_482_mask = 1'h1;
  assign mem_MPORT_482_en = reset;
  assign mem_MPORT_483_data = 19'h0;
  assign mem_MPORT_483_addr = 9'h1e3;
  assign mem_MPORT_483_mask = 1'h1;
  assign mem_MPORT_483_en = reset;
  assign mem_MPORT_484_data = 19'h0;
  assign mem_MPORT_484_addr = 9'h1e4;
  assign mem_MPORT_484_mask = 1'h1;
  assign mem_MPORT_484_en = reset;
  assign mem_MPORT_485_data = 19'h0;
  assign mem_MPORT_485_addr = 9'h1e5;
  assign mem_MPORT_485_mask = 1'h1;
  assign mem_MPORT_485_en = reset;
  assign mem_MPORT_486_data = 19'h0;
  assign mem_MPORT_486_addr = 9'h1e6;
  assign mem_MPORT_486_mask = 1'h1;
  assign mem_MPORT_486_en = reset;
  assign mem_MPORT_487_data = 19'h0;
  assign mem_MPORT_487_addr = 9'h1e7;
  assign mem_MPORT_487_mask = 1'h1;
  assign mem_MPORT_487_en = reset;
  assign mem_MPORT_488_data = 19'h0;
  assign mem_MPORT_488_addr = 9'h1e8;
  assign mem_MPORT_488_mask = 1'h1;
  assign mem_MPORT_488_en = reset;
  assign mem_MPORT_489_data = 19'h0;
  assign mem_MPORT_489_addr = 9'h1e9;
  assign mem_MPORT_489_mask = 1'h1;
  assign mem_MPORT_489_en = reset;
  assign mem_MPORT_490_data = 19'h0;
  assign mem_MPORT_490_addr = 9'h1ea;
  assign mem_MPORT_490_mask = 1'h1;
  assign mem_MPORT_490_en = reset;
  assign mem_MPORT_491_data = 19'h0;
  assign mem_MPORT_491_addr = 9'h1eb;
  assign mem_MPORT_491_mask = 1'h1;
  assign mem_MPORT_491_en = reset;
  assign mem_MPORT_492_data = 19'h0;
  assign mem_MPORT_492_addr = 9'h1ec;
  assign mem_MPORT_492_mask = 1'h1;
  assign mem_MPORT_492_en = reset;
  assign mem_MPORT_493_data = 19'h0;
  assign mem_MPORT_493_addr = 9'h1ed;
  assign mem_MPORT_493_mask = 1'h1;
  assign mem_MPORT_493_en = reset;
  assign mem_MPORT_494_data = 19'h0;
  assign mem_MPORT_494_addr = 9'h1ee;
  assign mem_MPORT_494_mask = 1'h1;
  assign mem_MPORT_494_en = reset;
  assign mem_MPORT_495_data = 19'h0;
  assign mem_MPORT_495_addr = 9'h1ef;
  assign mem_MPORT_495_mask = 1'h1;
  assign mem_MPORT_495_en = reset;
  assign mem_MPORT_496_data = 19'h0;
  assign mem_MPORT_496_addr = 9'h1f0;
  assign mem_MPORT_496_mask = 1'h1;
  assign mem_MPORT_496_en = reset;
  assign mem_MPORT_497_data = 19'h0;
  assign mem_MPORT_497_addr = 9'h1f1;
  assign mem_MPORT_497_mask = 1'h1;
  assign mem_MPORT_497_en = reset;
  assign mem_MPORT_498_data = 19'h0;
  assign mem_MPORT_498_addr = 9'h1f2;
  assign mem_MPORT_498_mask = 1'h1;
  assign mem_MPORT_498_en = reset;
  assign mem_MPORT_499_data = 19'h0;
  assign mem_MPORT_499_addr = 9'h1f3;
  assign mem_MPORT_499_mask = 1'h1;
  assign mem_MPORT_499_en = reset;
  assign mem_MPORT_500_data = 19'h0;
  assign mem_MPORT_500_addr = 9'h1f4;
  assign mem_MPORT_500_mask = 1'h1;
  assign mem_MPORT_500_en = reset;
  assign mem_MPORT_501_data = 19'h0;
  assign mem_MPORT_501_addr = 9'h1f5;
  assign mem_MPORT_501_mask = 1'h1;
  assign mem_MPORT_501_en = reset;
  assign mem_MPORT_502_data = 19'h0;
  assign mem_MPORT_502_addr = 9'h1f6;
  assign mem_MPORT_502_mask = 1'h1;
  assign mem_MPORT_502_en = reset;
  assign mem_MPORT_503_data = 19'h0;
  assign mem_MPORT_503_addr = 9'h1f7;
  assign mem_MPORT_503_mask = 1'h1;
  assign mem_MPORT_503_en = reset;
  assign mem_MPORT_504_data = 19'h0;
  assign mem_MPORT_504_addr = 9'h1f8;
  assign mem_MPORT_504_mask = 1'h1;
  assign mem_MPORT_504_en = reset;
  assign mem_MPORT_505_data = 19'h0;
  assign mem_MPORT_505_addr = 9'h1f9;
  assign mem_MPORT_505_mask = 1'h1;
  assign mem_MPORT_505_en = reset;
  assign mem_MPORT_506_data = 19'h0;
  assign mem_MPORT_506_addr = 9'h1fa;
  assign mem_MPORT_506_mask = 1'h1;
  assign mem_MPORT_506_en = reset;
  assign mem_MPORT_507_data = 19'h0;
  assign mem_MPORT_507_addr = 9'h1fb;
  assign mem_MPORT_507_mask = 1'h1;
  assign mem_MPORT_507_en = reset;
  assign mem_MPORT_508_data = 19'h0;
  assign mem_MPORT_508_addr = 9'h1fc;
  assign mem_MPORT_508_mask = 1'h1;
  assign mem_MPORT_508_en = reset;
  assign mem_MPORT_509_data = 19'h0;
  assign mem_MPORT_509_addr = 9'h1fd;
  assign mem_MPORT_509_mask = 1'h1;
  assign mem_MPORT_509_en = reset;
  assign mem_MPORT_510_data = 19'h0;
  assign mem_MPORT_510_addr = 9'h1fe;
  assign mem_MPORT_510_mask = 1'h1;
  assign mem_MPORT_510_en = reset;
  assign mem_MPORT_511_data = 19'h0;
  assign mem_MPORT_511_addr = 9'h1ff;
  assign mem_MPORT_511_mask = 1'h1;
  assign mem_MPORT_511_en = reset;
  assign mem_MPORT_512_data = io_w_data;
  assign mem_MPORT_512_addr = io_w_addr;
  assign mem_MPORT_512_mask = 1'h1;
  assign mem_MPORT_512_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_129_en & mem_MPORT_129_mask) begin
      mem[mem_MPORT_129_addr] <= mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_130_en & mem_MPORT_130_mask) begin
      mem[mem_MPORT_130_addr] <= mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_131_en & mem_MPORT_131_mask) begin
      mem[mem_MPORT_131_addr] <= mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_132_en & mem_MPORT_132_mask) begin
      mem[mem_MPORT_132_addr] <= mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_133_en & mem_MPORT_133_mask) begin
      mem[mem_MPORT_133_addr] <= mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_134_en & mem_MPORT_134_mask) begin
      mem[mem_MPORT_134_addr] <= mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_135_en & mem_MPORT_135_mask) begin
      mem[mem_MPORT_135_addr] <= mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_136_en & mem_MPORT_136_mask) begin
      mem[mem_MPORT_136_addr] <= mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_137_en & mem_MPORT_137_mask) begin
      mem[mem_MPORT_137_addr] <= mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_138_en & mem_MPORT_138_mask) begin
      mem[mem_MPORT_138_addr] <= mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_139_en & mem_MPORT_139_mask) begin
      mem[mem_MPORT_139_addr] <= mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_140_en & mem_MPORT_140_mask) begin
      mem[mem_MPORT_140_addr] <= mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_141_en & mem_MPORT_141_mask) begin
      mem[mem_MPORT_141_addr] <= mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_142_en & mem_MPORT_142_mask) begin
      mem[mem_MPORT_142_addr] <= mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_143_en & mem_MPORT_143_mask) begin
      mem[mem_MPORT_143_addr] <= mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_144_en & mem_MPORT_144_mask) begin
      mem[mem_MPORT_144_addr] <= mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_145_en & mem_MPORT_145_mask) begin
      mem[mem_MPORT_145_addr] <= mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_146_en & mem_MPORT_146_mask) begin
      mem[mem_MPORT_146_addr] <= mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_147_en & mem_MPORT_147_mask) begin
      mem[mem_MPORT_147_addr] <= mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_148_en & mem_MPORT_148_mask) begin
      mem[mem_MPORT_148_addr] <= mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_149_en & mem_MPORT_149_mask) begin
      mem[mem_MPORT_149_addr] <= mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_150_en & mem_MPORT_150_mask) begin
      mem[mem_MPORT_150_addr] <= mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_151_en & mem_MPORT_151_mask) begin
      mem[mem_MPORT_151_addr] <= mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_152_en & mem_MPORT_152_mask) begin
      mem[mem_MPORT_152_addr] <= mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_153_en & mem_MPORT_153_mask) begin
      mem[mem_MPORT_153_addr] <= mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_154_en & mem_MPORT_154_mask) begin
      mem[mem_MPORT_154_addr] <= mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_155_en & mem_MPORT_155_mask) begin
      mem[mem_MPORT_155_addr] <= mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_156_en & mem_MPORT_156_mask) begin
      mem[mem_MPORT_156_addr] <= mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_157_en & mem_MPORT_157_mask) begin
      mem[mem_MPORT_157_addr] <= mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_158_en & mem_MPORT_158_mask) begin
      mem[mem_MPORT_158_addr] <= mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_159_en & mem_MPORT_159_mask) begin
      mem[mem_MPORT_159_addr] <= mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_160_en & mem_MPORT_160_mask) begin
      mem[mem_MPORT_160_addr] <= mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_161_en & mem_MPORT_161_mask) begin
      mem[mem_MPORT_161_addr] <= mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_162_en & mem_MPORT_162_mask) begin
      mem[mem_MPORT_162_addr] <= mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_163_en & mem_MPORT_163_mask) begin
      mem[mem_MPORT_163_addr] <= mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_164_en & mem_MPORT_164_mask) begin
      mem[mem_MPORT_164_addr] <= mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_165_en & mem_MPORT_165_mask) begin
      mem[mem_MPORT_165_addr] <= mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_166_en & mem_MPORT_166_mask) begin
      mem[mem_MPORT_166_addr] <= mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_167_en & mem_MPORT_167_mask) begin
      mem[mem_MPORT_167_addr] <= mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_168_en & mem_MPORT_168_mask) begin
      mem[mem_MPORT_168_addr] <= mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_169_en & mem_MPORT_169_mask) begin
      mem[mem_MPORT_169_addr] <= mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_170_en & mem_MPORT_170_mask) begin
      mem[mem_MPORT_170_addr] <= mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_171_en & mem_MPORT_171_mask) begin
      mem[mem_MPORT_171_addr] <= mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_172_en & mem_MPORT_172_mask) begin
      mem[mem_MPORT_172_addr] <= mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_173_en & mem_MPORT_173_mask) begin
      mem[mem_MPORT_173_addr] <= mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_174_en & mem_MPORT_174_mask) begin
      mem[mem_MPORT_174_addr] <= mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_175_en & mem_MPORT_175_mask) begin
      mem[mem_MPORT_175_addr] <= mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_176_en & mem_MPORT_176_mask) begin
      mem[mem_MPORT_176_addr] <= mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_177_en & mem_MPORT_177_mask) begin
      mem[mem_MPORT_177_addr] <= mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_178_en & mem_MPORT_178_mask) begin
      mem[mem_MPORT_178_addr] <= mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_179_en & mem_MPORT_179_mask) begin
      mem[mem_MPORT_179_addr] <= mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_180_en & mem_MPORT_180_mask) begin
      mem[mem_MPORT_180_addr] <= mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_181_en & mem_MPORT_181_mask) begin
      mem[mem_MPORT_181_addr] <= mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_182_en & mem_MPORT_182_mask) begin
      mem[mem_MPORT_182_addr] <= mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_183_en & mem_MPORT_183_mask) begin
      mem[mem_MPORT_183_addr] <= mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_184_en & mem_MPORT_184_mask) begin
      mem[mem_MPORT_184_addr] <= mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_185_en & mem_MPORT_185_mask) begin
      mem[mem_MPORT_185_addr] <= mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_186_en & mem_MPORT_186_mask) begin
      mem[mem_MPORT_186_addr] <= mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_187_en & mem_MPORT_187_mask) begin
      mem[mem_MPORT_187_addr] <= mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_188_en & mem_MPORT_188_mask) begin
      mem[mem_MPORT_188_addr] <= mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_189_en & mem_MPORT_189_mask) begin
      mem[mem_MPORT_189_addr] <= mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_190_en & mem_MPORT_190_mask) begin
      mem[mem_MPORT_190_addr] <= mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_191_en & mem_MPORT_191_mask) begin
      mem[mem_MPORT_191_addr] <= mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_192_en & mem_MPORT_192_mask) begin
      mem[mem_MPORT_192_addr] <= mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_193_en & mem_MPORT_193_mask) begin
      mem[mem_MPORT_193_addr] <= mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_194_en & mem_MPORT_194_mask) begin
      mem[mem_MPORT_194_addr] <= mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_195_en & mem_MPORT_195_mask) begin
      mem[mem_MPORT_195_addr] <= mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_196_en & mem_MPORT_196_mask) begin
      mem[mem_MPORT_196_addr] <= mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_197_en & mem_MPORT_197_mask) begin
      mem[mem_MPORT_197_addr] <= mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_198_en & mem_MPORT_198_mask) begin
      mem[mem_MPORT_198_addr] <= mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_199_en & mem_MPORT_199_mask) begin
      mem[mem_MPORT_199_addr] <= mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_200_en & mem_MPORT_200_mask) begin
      mem[mem_MPORT_200_addr] <= mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_201_en & mem_MPORT_201_mask) begin
      mem[mem_MPORT_201_addr] <= mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_202_en & mem_MPORT_202_mask) begin
      mem[mem_MPORT_202_addr] <= mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_203_en & mem_MPORT_203_mask) begin
      mem[mem_MPORT_203_addr] <= mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_204_en & mem_MPORT_204_mask) begin
      mem[mem_MPORT_204_addr] <= mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_205_en & mem_MPORT_205_mask) begin
      mem[mem_MPORT_205_addr] <= mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_206_en & mem_MPORT_206_mask) begin
      mem[mem_MPORT_206_addr] <= mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_207_en & mem_MPORT_207_mask) begin
      mem[mem_MPORT_207_addr] <= mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_208_en & mem_MPORT_208_mask) begin
      mem[mem_MPORT_208_addr] <= mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_209_en & mem_MPORT_209_mask) begin
      mem[mem_MPORT_209_addr] <= mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_210_en & mem_MPORT_210_mask) begin
      mem[mem_MPORT_210_addr] <= mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_211_en & mem_MPORT_211_mask) begin
      mem[mem_MPORT_211_addr] <= mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_212_en & mem_MPORT_212_mask) begin
      mem[mem_MPORT_212_addr] <= mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_213_en & mem_MPORT_213_mask) begin
      mem[mem_MPORT_213_addr] <= mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_214_en & mem_MPORT_214_mask) begin
      mem[mem_MPORT_214_addr] <= mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_215_en & mem_MPORT_215_mask) begin
      mem[mem_MPORT_215_addr] <= mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_216_en & mem_MPORT_216_mask) begin
      mem[mem_MPORT_216_addr] <= mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_217_en & mem_MPORT_217_mask) begin
      mem[mem_MPORT_217_addr] <= mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_218_en & mem_MPORT_218_mask) begin
      mem[mem_MPORT_218_addr] <= mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_219_en & mem_MPORT_219_mask) begin
      mem[mem_MPORT_219_addr] <= mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_220_en & mem_MPORT_220_mask) begin
      mem[mem_MPORT_220_addr] <= mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_221_en & mem_MPORT_221_mask) begin
      mem[mem_MPORT_221_addr] <= mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_222_en & mem_MPORT_222_mask) begin
      mem[mem_MPORT_222_addr] <= mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_223_en & mem_MPORT_223_mask) begin
      mem[mem_MPORT_223_addr] <= mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_224_en & mem_MPORT_224_mask) begin
      mem[mem_MPORT_224_addr] <= mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_225_en & mem_MPORT_225_mask) begin
      mem[mem_MPORT_225_addr] <= mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_226_en & mem_MPORT_226_mask) begin
      mem[mem_MPORT_226_addr] <= mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_227_en & mem_MPORT_227_mask) begin
      mem[mem_MPORT_227_addr] <= mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_228_en & mem_MPORT_228_mask) begin
      mem[mem_MPORT_228_addr] <= mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_229_en & mem_MPORT_229_mask) begin
      mem[mem_MPORT_229_addr] <= mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_230_en & mem_MPORT_230_mask) begin
      mem[mem_MPORT_230_addr] <= mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_231_en & mem_MPORT_231_mask) begin
      mem[mem_MPORT_231_addr] <= mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_232_en & mem_MPORT_232_mask) begin
      mem[mem_MPORT_232_addr] <= mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_233_en & mem_MPORT_233_mask) begin
      mem[mem_MPORT_233_addr] <= mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_234_en & mem_MPORT_234_mask) begin
      mem[mem_MPORT_234_addr] <= mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_235_en & mem_MPORT_235_mask) begin
      mem[mem_MPORT_235_addr] <= mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_236_en & mem_MPORT_236_mask) begin
      mem[mem_MPORT_236_addr] <= mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_237_en & mem_MPORT_237_mask) begin
      mem[mem_MPORT_237_addr] <= mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_238_en & mem_MPORT_238_mask) begin
      mem[mem_MPORT_238_addr] <= mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_239_en & mem_MPORT_239_mask) begin
      mem[mem_MPORT_239_addr] <= mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_240_en & mem_MPORT_240_mask) begin
      mem[mem_MPORT_240_addr] <= mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_241_en & mem_MPORT_241_mask) begin
      mem[mem_MPORT_241_addr] <= mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_242_en & mem_MPORT_242_mask) begin
      mem[mem_MPORT_242_addr] <= mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_243_en & mem_MPORT_243_mask) begin
      mem[mem_MPORT_243_addr] <= mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_244_en & mem_MPORT_244_mask) begin
      mem[mem_MPORT_244_addr] <= mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_245_en & mem_MPORT_245_mask) begin
      mem[mem_MPORT_245_addr] <= mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_246_en & mem_MPORT_246_mask) begin
      mem[mem_MPORT_246_addr] <= mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_247_en & mem_MPORT_247_mask) begin
      mem[mem_MPORT_247_addr] <= mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_248_en & mem_MPORT_248_mask) begin
      mem[mem_MPORT_248_addr] <= mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_249_en & mem_MPORT_249_mask) begin
      mem[mem_MPORT_249_addr] <= mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_250_en & mem_MPORT_250_mask) begin
      mem[mem_MPORT_250_addr] <= mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_251_en & mem_MPORT_251_mask) begin
      mem[mem_MPORT_251_addr] <= mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_252_en & mem_MPORT_252_mask) begin
      mem[mem_MPORT_252_addr] <= mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_253_en & mem_MPORT_253_mask) begin
      mem[mem_MPORT_253_addr] <= mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_254_en & mem_MPORT_254_mask) begin
      mem[mem_MPORT_254_addr] <= mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_255_en & mem_MPORT_255_mask) begin
      mem[mem_MPORT_255_addr] <= mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_256_en & mem_MPORT_256_mask) begin
      mem[mem_MPORT_256_addr] <= mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_257_en & mem_MPORT_257_mask) begin
      mem[mem_MPORT_257_addr] <= mem_MPORT_257_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_258_en & mem_MPORT_258_mask) begin
      mem[mem_MPORT_258_addr] <= mem_MPORT_258_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_259_en & mem_MPORT_259_mask) begin
      mem[mem_MPORT_259_addr] <= mem_MPORT_259_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_260_en & mem_MPORT_260_mask) begin
      mem[mem_MPORT_260_addr] <= mem_MPORT_260_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_261_en & mem_MPORT_261_mask) begin
      mem[mem_MPORT_261_addr] <= mem_MPORT_261_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_262_en & mem_MPORT_262_mask) begin
      mem[mem_MPORT_262_addr] <= mem_MPORT_262_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_263_en & mem_MPORT_263_mask) begin
      mem[mem_MPORT_263_addr] <= mem_MPORT_263_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_264_en & mem_MPORT_264_mask) begin
      mem[mem_MPORT_264_addr] <= mem_MPORT_264_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_265_en & mem_MPORT_265_mask) begin
      mem[mem_MPORT_265_addr] <= mem_MPORT_265_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_266_en & mem_MPORT_266_mask) begin
      mem[mem_MPORT_266_addr] <= mem_MPORT_266_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_267_en & mem_MPORT_267_mask) begin
      mem[mem_MPORT_267_addr] <= mem_MPORT_267_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_268_en & mem_MPORT_268_mask) begin
      mem[mem_MPORT_268_addr] <= mem_MPORT_268_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_269_en & mem_MPORT_269_mask) begin
      mem[mem_MPORT_269_addr] <= mem_MPORT_269_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_270_en & mem_MPORT_270_mask) begin
      mem[mem_MPORT_270_addr] <= mem_MPORT_270_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_271_en & mem_MPORT_271_mask) begin
      mem[mem_MPORT_271_addr] <= mem_MPORT_271_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_272_en & mem_MPORT_272_mask) begin
      mem[mem_MPORT_272_addr] <= mem_MPORT_272_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_273_en & mem_MPORT_273_mask) begin
      mem[mem_MPORT_273_addr] <= mem_MPORT_273_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_274_en & mem_MPORT_274_mask) begin
      mem[mem_MPORT_274_addr] <= mem_MPORT_274_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_275_en & mem_MPORT_275_mask) begin
      mem[mem_MPORT_275_addr] <= mem_MPORT_275_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_276_en & mem_MPORT_276_mask) begin
      mem[mem_MPORT_276_addr] <= mem_MPORT_276_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_277_en & mem_MPORT_277_mask) begin
      mem[mem_MPORT_277_addr] <= mem_MPORT_277_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_278_en & mem_MPORT_278_mask) begin
      mem[mem_MPORT_278_addr] <= mem_MPORT_278_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_279_en & mem_MPORT_279_mask) begin
      mem[mem_MPORT_279_addr] <= mem_MPORT_279_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_280_en & mem_MPORT_280_mask) begin
      mem[mem_MPORT_280_addr] <= mem_MPORT_280_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_281_en & mem_MPORT_281_mask) begin
      mem[mem_MPORT_281_addr] <= mem_MPORT_281_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_282_en & mem_MPORT_282_mask) begin
      mem[mem_MPORT_282_addr] <= mem_MPORT_282_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_283_en & mem_MPORT_283_mask) begin
      mem[mem_MPORT_283_addr] <= mem_MPORT_283_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_284_en & mem_MPORT_284_mask) begin
      mem[mem_MPORT_284_addr] <= mem_MPORT_284_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_285_en & mem_MPORT_285_mask) begin
      mem[mem_MPORT_285_addr] <= mem_MPORT_285_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_286_en & mem_MPORT_286_mask) begin
      mem[mem_MPORT_286_addr] <= mem_MPORT_286_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_287_en & mem_MPORT_287_mask) begin
      mem[mem_MPORT_287_addr] <= mem_MPORT_287_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_288_en & mem_MPORT_288_mask) begin
      mem[mem_MPORT_288_addr] <= mem_MPORT_288_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_289_en & mem_MPORT_289_mask) begin
      mem[mem_MPORT_289_addr] <= mem_MPORT_289_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_290_en & mem_MPORT_290_mask) begin
      mem[mem_MPORT_290_addr] <= mem_MPORT_290_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_291_en & mem_MPORT_291_mask) begin
      mem[mem_MPORT_291_addr] <= mem_MPORT_291_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_292_en & mem_MPORT_292_mask) begin
      mem[mem_MPORT_292_addr] <= mem_MPORT_292_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_293_en & mem_MPORT_293_mask) begin
      mem[mem_MPORT_293_addr] <= mem_MPORT_293_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_294_en & mem_MPORT_294_mask) begin
      mem[mem_MPORT_294_addr] <= mem_MPORT_294_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_295_en & mem_MPORT_295_mask) begin
      mem[mem_MPORT_295_addr] <= mem_MPORT_295_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_296_en & mem_MPORT_296_mask) begin
      mem[mem_MPORT_296_addr] <= mem_MPORT_296_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_297_en & mem_MPORT_297_mask) begin
      mem[mem_MPORT_297_addr] <= mem_MPORT_297_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_298_en & mem_MPORT_298_mask) begin
      mem[mem_MPORT_298_addr] <= mem_MPORT_298_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_299_en & mem_MPORT_299_mask) begin
      mem[mem_MPORT_299_addr] <= mem_MPORT_299_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_300_en & mem_MPORT_300_mask) begin
      mem[mem_MPORT_300_addr] <= mem_MPORT_300_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_301_en & mem_MPORT_301_mask) begin
      mem[mem_MPORT_301_addr] <= mem_MPORT_301_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_302_en & mem_MPORT_302_mask) begin
      mem[mem_MPORT_302_addr] <= mem_MPORT_302_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_303_en & mem_MPORT_303_mask) begin
      mem[mem_MPORT_303_addr] <= mem_MPORT_303_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_304_en & mem_MPORT_304_mask) begin
      mem[mem_MPORT_304_addr] <= mem_MPORT_304_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_305_en & mem_MPORT_305_mask) begin
      mem[mem_MPORT_305_addr] <= mem_MPORT_305_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_306_en & mem_MPORT_306_mask) begin
      mem[mem_MPORT_306_addr] <= mem_MPORT_306_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_307_en & mem_MPORT_307_mask) begin
      mem[mem_MPORT_307_addr] <= mem_MPORT_307_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_308_en & mem_MPORT_308_mask) begin
      mem[mem_MPORT_308_addr] <= mem_MPORT_308_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_309_en & mem_MPORT_309_mask) begin
      mem[mem_MPORT_309_addr] <= mem_MPORT_309_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_310_en & mem_MPORT_310_mask) begin
      mem[mem_MPORT_310_addr] <= mem_MPORT_310_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_311_en & mem_MPORT_311_mask) begin
      mem[mem_MPORT_311_addr] <= mem_MPORT_311_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_312_en & mem_MPORT_312_mask) begin
      mem[mem_MPORT_312_addr] <= mem_MPORT_312_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_313_en & mem_MPORT_313_mask) begin
      mem[mem_MPORT_313_addr] <= mem_MPORT_313_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_314_en & mem_MPORT_314_mask) begin
      mem[mem_MPORT_314_addr] <= mem_MPORT_314_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_315_en & mem_MPORT_315_mask) begin
      mem[mem_MPORT_315_addr] <= mem_MPORT_315_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_316_en & mem_MPORT_316_mask) begin
      mem[mem_MPORT_316_addr] <= mem_MPORT_316_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_317_en & mem_MPORT_317_mask) begin
      mem[mem_MPORT_317_addr] <= mem_MPORT_317_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_318_en & mem_MPORT_318_mask) begin
      mem[mem_MPORT_318_addr] <= mem_MPORT_318_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_319_en & mem_MPORT_319_mask) begin
      mem[mem_MPORT_319_addr] <= mem_MPORT_319_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_320_en & mem_MPORT_320_mask) begin
      mem[mem_MPORT_320_addr] <= mem_MPORT_320_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_321_en & mem_MPORT_321_mask) begin
      mem[mem_MPORT_321_addr] <= mem_MPORT_321_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_322_en & mem_MPORT_322_mask) begin
      mem[mem_MPORT_322_addr] <= mem_MPORT_322_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_323_en & mem_MPORT_323_mask) begin
      mem[mem_MPORT_323_addr] <= mem_MPORT_323_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_324_en & mem_MPORT_324_mask) begin
      mem[mem_MPORT_324_addr] <= mem_MPORT_324_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_325_en & mem_MPORT_325_mask) begin
      mem[mem_MPORT_325_addr] <= mem_MPORT_325_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_326_en & mem_MPORT_326_mask) begin
      mem[mem_MPORT_326_addr] <= mem_MPORT_326_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_327_en & mem_MPORT_327_mask) begin
      mem[mem_MPORT_327_addr] <= mem_MPORT_327_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_328_en & mem_MPORT_328_mask) begin
      mem[mem_MPORT_328_addr] <= mem_MPORT_328_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_329_en & mem_MPORT_329_mask) begin
      mem[mem_MPORT_329_addr] <= mem_MPORT_329_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_330_en & mem_MPORT_330_mask) begin
      mem[mem_MPORT_330_addr] <= mem_MPORT_330_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_331_en & mem_MPORT_331_mask) begin
      mem[mem_MPORT_331_addr] <= mem_MPORT_331_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_332_en & mem_MPORT_332_mask) begin
      mem[mem_MPORT_332_addr] <= mem_MPORT_332_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_333_en & mem_MPORT_333_mask) begin
      mem[mem_MPORT_333_addr] <= mem_MPORT_333_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_334_en & mem_MPORT_334_mask) begin
      mem[mem_MPORT_334_addr] <= mem_MPORT_334_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_335_en & mem_MPORT_335_mask) begin
      mem[mem_MPORT_335_addr] <= mem_MPORT_335_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_336_en & mem_MPORT_336_mask) begin
      mem[mem_MPORT_336_addr] <= mem_MPORT_336_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_337_en & mem_MPORT_337_mask) begin
      mem[mem_MPORT_337_addr] <= mem_MPORT_337_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_338_en & mem_MPORT_338_mask) begin
      mem[mem_MPORT_338_addr] <= mem_MPORT_338_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_339_en & mem_MPORT_339_mask) begin
      mem[mem_MPORT_339_addr] <= mem_MPORT_339_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_340_en & mem_MPORT_340_mask) begin
      mem[mem_MPORT_340_addr] <= mem_MPORT_340_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_341_en & mem_MPORT_341_mask) begin
      mem[mem_MPORT_341_addr] <= mem_MPORT_341_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_342_en & mem_MPORT_342_mask) begin
      mem[mem_MPORT_342_addr] <= mem_MPORT_342_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_343_en & mem_MPORT_343_mask) begin
      mem[mem_MPORT_343_addr] <= mem_MPORT_343_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_344_en & mem_MPORT_344_mask) begin
      mem[mem_MPORT_344_addr] <= mem_MPORT_344_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_345_en & mem_MPORT_345_mask) begin
      mem[mem_MPORT_345_addr] <= mem_MPORT_345_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_346_en & mem_MPORT_346_mask) begin
      mem[mem_MPORT_346_addr] <= mem_MPORT_346_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_347_en & mem_MPORT_347_mask) begin
      mem[mem_MPORT_347_addr] <= mem_MPORT_347_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_348_en & mem_MPORT_348_mask) begin
      mem[mem_MPORT_348_addr] <= mem_MPORT_348_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_349_en & mem_MPORT_349_mask) begin
      mem[mem_MPORT_349_addr] <= mem_MPORT_349_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_350_en & mem_MPORT_350_mask) begin
      mem[mem_MPORT_350_addr] <= mem_MPORT_350_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_351_en & mem_MPORT_351_mask) begin
      mem[mem_MPORT_351_addr] <= mem_MPORT_351_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_352_en & mem_MPORT_352_mask) begin
      mem[mem_MPORT_352_addr] <= mem_MPORT_352_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_353_en & mem_MPORT_353_mask) begin
      mem[mem_MPORT_353_addr] <= mem_MPORT_353_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_354_en & mem_MPORT_354_mask) begin
      mem[mem_MPORT_354_addr] <= mem_MPORT_354_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_355_en & mem_MPORT_355_mask) begin
      mem[mem_MPORT_355_addr] <= mem_MPORT_355_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_356_en & mem_MPORT_356_mask) begin
      mem[mem_MPORT_356_addr] <= mem_MPORT_356_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_357_en & mem_MPORT_357_mask) begin
      mem[mem_MPORT_357_addr] <= mem_MPORT_357_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_358_en & mem_MPORT_358_mask) begin
      mem[mem_MPORT_358_addr] <= mem_MPORT_358_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_359_en & mem_MPORT_359_mask) begin
      mem[mem_MPORT_359_addr] <= mem_MPORT_359_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_360_en & mem_MPORT_360_mask) begin
      mem[mem_MPORT_360_addr] <= mem_MPORT_360_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_361_en & mem_MPORT_361_mask) begin
      mem[mem_MPORT_361_addr] <= mem_MPORT_361_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_362_en & mem_MPORT_362_mask) begin
      mem[mem_MPORT_362_addr] <= mem_MPORT_362_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_363_en & mem_MPORT_363_mask) begin
      mem[mem_MPORT_363_addr] <= mem_MPORT_363_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_364_en & mem_MPORT_364_mask) begin
      mem[mem_MPORT_364_addr] <= mem_MPORT_364_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_365_en & mem_MPORT_365_mask) begin
      mem[mem_MPORT_365_addr] <= mem_MPORT_365_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_366_en & mem_MPORT_366_mask) begin
      mem[mem_MPORT_366_addr] <= mem_MPORT_366_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_367_en & mem_MPORT_367_mask) begin
      mem[mem_MPORT_367_addr] <= mem_MPORT_367_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_368_en & mem_MPORT_368_mask) begin
      mem[mem_MPORT_368_addr] <= mem_MPORT_368_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_369_en & mem_MPORT_369_mask) begin
      mem[mem_MPORT_369_addr] <= mem_MPORT_369_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_370_en & mem_MPORT_370_mask) begin
      mem[mem_MPORT_370_addr] <= mem_MPORT_370_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_371_en & mem_MPORT_371_mask) begin
      mem[mem_MPORT_371_addr] <= mem_MPORT_371_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_372_en & mem_MPORT_372_mask) begin
      mem[mem_MPORT_372_addr] <= mem_MPORT_372_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_373_en & mem_MPORT_373_mask) begin
      mem[mem_MPORT_373_addr] <= mem_MPORT_373_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_374_en & mem_MPORT_374_mask) begin
      mem[mem_MPORT_374_addr] <= mem_MPORT_374_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_375_en & mem_MPORT_375_mask) begin
      mem[mem_MPORT_375_addr] <= mem_MPORT_375_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_376_en & mem_MPORT_376_mask) begin
      mem[mem_MPORT_376_addr] <= mem_MPORT_376_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_377_en & mem_MPORT_377_mask) begin
      mem[mem_MPORT_377_addr] <= mem_MPORT_377_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_378_en & mem_MPORT_378_mask) begin
      mem[mem_MPORT_378_addr] <= mem_MPORT_378_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_379_en & mem_MPORT_379_mask) begin
      mem[mem_MPORT_379_addr] <= mem_MPORT_379_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_380_en & mem_MPORT_380_mask) begin
      mem[mem_MPORT_380_addr] <= mem_MPORT_380_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_381_en & mem_MPORT_381_mask) begin
      mem[mem_MPORT_381_addr] <= mem_MPORT_381_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_382_en & mem_MPORT_382_mask) begin
      mem[mem_MPORT_382_addr] <= mem_MPORT_382_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_383_en & mem_MPORT_383_mask) begin
      mem[mem_MPORT_383_addr] <= mem_MPORT_383_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_384_en & mem_MPORT_384_mask) begin
      mem[mem_MPORT_384_addr] <= mem_MPORT_384_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_385_en & mem_MPORT_385_mask) begin
      mem[mem_MPORT_385_addr] <= mem_MPORT_385_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_386_en & mem_MPORT_386_mask) begin
      mem[mem_MPORT_386_addr] <= mem_MPORT_386_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_387_en & mem_MPORT_387_mask) begin
      mem[mem_MPORT_387_addr] <= mem_MPORT_387_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_388_en & mem_MPORT_388_mask) begin
      mem[mem_MPORT_388_addr] <= mem_MPORT_388_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_389_en & mem_MPORT_389_mask) begin
      mem[mem_MPORT_389_addr] <= mem_MPORT_389_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_390_en & mem_MPORT_390_mask) begin
      mem[mem_MPORT_390_addr] <= mem_MPORT_390_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_391_en & mem_MPORT_391_mask) begin
      mem[mem_MPORT_391_addr] <= mem_MPORT_391_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_392_en & mem_MPORT_392_mask) begin
      mem[mem_MPORT_392_addr] <= mem_MPORT_392_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_393_en & mem_MPORT_393_mask) begin
      mem[mem_MPORT_393_addr] <= mem_MPORT_393_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_394_en & mem_MPORT_394_mask) begin
      mem[mem_MPORT_394_addr] <= mem_MPORT_394_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_395_en & mem_MPORT_395_mask) begin
      mem[mem_MPORT_395_addr] <= mem_MPORT_395_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_396_en & mem_MPORT_396_mask) begin
      mem[mem_MPORT_396_addr] <= mem_MPORT_396_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_397_en & mem_MPORT_397_mask) begin
      mem[mem_MPORT_397_addr] <= mem_MPORT_397_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_398_en & mem_MPORT_398_mask) begin
      mem[mem_MPORT_398_addr] <= mem_MPORT_398_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_399_en & mem_MPORT_399_mask) begin
      mem[mem_MPORT_399_addr] <= mem_MPORT_399_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_400_en & mem_MPORT_400_mask) begin
      mem[mem_MPORT_400_addr] <= mem_MPORT_400_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_401_en & mem_MPORT_401_mask) begin
      mem[mem_MPORT_401_addr] <= mem_MPORT_401_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_402_en & mem_MPORT_402_mask) begin
      mem[mem_MPORT_402_addr] <= mem_MPORT_402_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_403_en & mem_MPORT_403_mask) begin
      mem[mem_MPORT_403_addr] <= mem_MPORT_403_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_404_en & mem_MPORT_404_mask) begin
      mem[mem_MPORT_404_addr] <= mem_MPORT_404_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_405_en & mem_MPORT_405_mask) begin
      mem[mem_MPORT_405_addr] <= mem_MPORT_405_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_406_en & mem_MPORT_406_mask) begin
      mem[mem_MPORT_406_addr] <= mem_MPORT_406_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_407_en & mem_MPORT_407_mask) begin
      mem[mem_MPORT_407_addr] <= mem_MPORT_407_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_408_en & mem_MPORT_408_mask) begin
      mem[mem_MPORT_408_addr] <= mem_MPORT_408_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_409_en & mem_MPORT_409_mask) begin
      mem[mem_MPORT_409_addr] <= mem_MPORT_409_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_410_en & mem_MPORT_410_mask) begin
      mem[mem_MPORT_410_addr] <= mem_MPORT_410_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_411_en & mem_MPORT_411_mask) begin
      mem[mem_MPORT_411_addr] <= mem_MPORT_411_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_412_en & mem_MPORT_412_mask) begin
      mem[mem_MPORT_412_addr] <= mem_MPORT_412_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_413_en & mem_MPORT_413_mask) begin
      mem[mem_MPORT_413_addr] <= mem_MPORT_413_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_414_en & mem_MPORT_414_mask) begin
      mem[mem_MPORT_414_addr] <= mem_MPORT_414_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_415_en & mem_MPORT_415_mask) begin
      mem[mem_MPORT_415_addr] <= mem_MPORT_415_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_416_en & mem_MPORT_416_mask) begin
      mem[mem_MPORT_416_addr] <= mem_MPORT_416_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_417_en & mem_MPORT_417_mask) begin
      mem[mem_MPORT_417_addr] <= mem_MPORT_417_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_418_en & mem_MPORT_418_mask) begin
      mem[mem_MPORT_418_addr] <= mem_MPORT_418_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_419_en & mem_MPORT_419_mask) begin
      mem[mem_MPORT_419_addr] <= mem_MPORT_419_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_420_en & mem_MPORT_420_mask) begin
      mem[mem_MPORT_420_addr] <= mem_MPORT_420_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_421_en & mem_MPORT_421_mask) begin
      mem[mem_MPORT_421_addr] <= mem_MPORT_421_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_422_en & mem_MPORT_422_mask) begin
      mem[mem_MPORT_422_addr] <= mem_MPORT_422_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_423_en & mem_MPORT_423_mask) begin
      mem[mem_MPORT_423_addr] <= mem_MPORT_423_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_424_en & mem_MPORT_424_mask) begin
      mem[mem_MPORT_424_addr] <= mem_MPORT_424_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_425_en & mem_MPORT_425_mask) begin
      mem[mem_MPORT_425_addr] <= mem_MPORT_425_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_426_en & mem_MPORT_426_mask) begin
      mem[mem_MPORT_426_addr] <= mem_MPORT_426_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_427_en & mem_MPORT_427_mask) begin
      mem[mem_MPORT_427_addr] <= mem_MPORT_427_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_428_en & mem_MPORT_428_mask) begin
      mem[mem_MPORT_428_addr] <= mem_MPORT_428_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_429_en & mem_MPORT_429_mask) begin
      mem[mem_MPORT_429_addr] <= mem_MPORT_429_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_430_en & mem_MPORT_430_mask) begin
      mem[mem_MPORT_430_addr] <= mem_MPORT_430_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_431_en & mem_MPORT_431_mask) begin
      mem[mem_MPORT_431_addr] <= mem_MPORT_431_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_432_en & mem_MPORT_432_mask) begin
      mem[mem_MPORT_432_addr] <= mem_MPORT_432_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_433_en & mem_MPORT_433_mask) begin
      mem[mem_MPORT_433_addr] <= mem_MPORT_433_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_434_en & mem_MPORT_434_mask) begin
      mem[mem_MPORT_434_addr] <= mem_MPORT_434_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_435_en & mem_MPORT_435_mask) begin
      mem[mem_MPORT_435_addr] <= mem_MPORT_435_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_436_en & mem_MPORT_436_mask) begin
      mem[mem_MPORT_436_addr] <= mem_MPORT_436_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_437_en & mem_MPORT_437_mask) begin
      mem[mem_MPORT_437_addr] <= mem_MPORT_437_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_438_en & mem_MPORT_438_mask) begin
      mem[mem_MPORT_438_addr] <= mem_MPORT_438_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_439_en & mem_MPORT_439_mask) begin
      mem[mem_MPORT_439_addr] <= mem_MPORT_439_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_440_en & mem_MPORT_440_mask) begin
      mem[mem_MPORT_440_addr] <= mem_MPORT_440_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_441_en & mem_MPORT_441_mask) begin
      mem[mem_MPORT_441_addr] <= mem_MPORT_441_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_442_en & mem_MPORT_442_mask) begin
      mem[mem_MPORT_442_addr] <= mem_MPORT_442_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_443_en & mem_MPORT_443_mask) begin
      mem[mem_MPORT_443_addr] <= mem_MPORT_443_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_444_en & mem_MPORT_444_mask) begin
      mem[mem_MPORT_444_addr] <= mem_MPORT_444_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_445_en & mem_MPORT_445_mask) begin
      mem[mem_MPORT_445_addr] <= mem_MPORT_445_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_446_en & mem_MPORT_446_mask) begin
      mem[mem_MPORT_446_addr] <= mem_MPORT_446_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_447_en & mem_MPORT_447_mask) begin
      mem[mem_MPORT_447_addr] <= mem_MPORT_447_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_448_en & mem_MPORT_448_mask) begin
      mem[mem_MPORT_448_addr] <= mem_MPORT_448_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_449_en & mem_MPORT_449_mask) begin
      mem[mem_MPORT_449_addr] <= mem_MPORT_449_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_450_en & mem_MPORT_450_mask) begin
      mem[mem_MPORT_450_addr] <= mem_MPORT_450_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_451_en & mem_MPORT_451_mask) begin
      mem[mem_MPORT_451_addr] <= mem_MPORT_451_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_452_en & mem_MPORT_452_mask) begin
      mem[mem_MPORT_452_addr] <= mem_MPORT_452_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_453_en & mem_MPORT_453_mask) begin
      mem[mem_MPORT_453_addr] <= mem_MPORT_453_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_454_en & mem_MPORT_454_mask) begin
      mem[mem_MPORT_454_addr] <= mem_MPORT_454_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_455_en & mem_MPORT_455_mask) begin
      mem[mem_MPORT_455_addr] <= mem_MPORT_455_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_456_en & mem_MPORT_456_mask) begin
      mem[mem_MPORT_456_addr] <= mem_MPORT_456_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_457_en & mem_MPORT_457_mask) begin
      mem[mem_MPORT_457_addr] <= mem_MPORT_457_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_458_en & mem_MPORT_458_mask) begin
      mem[mem_MPORT_458_addr] <= mem_MPORT_458_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_459_en & mem_MPORT_459_mask) begin
      mem[mem_MPORT_459_addr] <= mem_MPORT_459_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_460_en & mem_MPORT_460_mask) begin
      mem[mem_MPORT_460_addr] <= mem_MPORT_460_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_461_en & mem_MPORT_461_mask) begin
      mem[mem_MPORT_461_addr] <= mem_MPORT_461_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_462_en & mem_MPORT_462_mask) begin
      mem[mem_MPORT_462_addr] <= mem_MPORT_462_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_463_en & mem_MPORT_463_mask) begin
      mem[mem_MPORT_463_addr] <= mem_MPORT_463_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_464_en & mem_MPORT_464_mask) begin
      mem[mem_MPORT_464_addr] <= mem_MPORT_464_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_465_en & mem_MPORT_465_mask) begin
      mem[mem_MPORT_465_addr] <= mem_MPORT_465_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_466_en & mem_MPORT_466_mask) begin
      mem[mem_MPORT_466_addr] <= mem_MPORT_466_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_467_en & mem_MPORT_467_mask) begin
      mem[mem_MPORT_467_addr] <= mem_MPORT_467_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_468_en & mem_MPORT_468_mask) begin
      mem[mem_MPORT_468_addr] <= mem_MPORT_468_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_469_en & mem_MPORT_469_mask) begin
      mem[mem_MPORT_469_addr] <= mem_MPORT_469_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_470_en & mem_MPORT_470_mask) begin
      mem[mem_MPORT_470_addr] <= mem_MPORT_470_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_471_en & mem_MPORT_471_mask) begin
      mem[mem_MPORT_471_addr] <= mem_MPORT_471_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_472_en & mem_MPORT_472_mask) begin
      mem[mem_MPORT_472_addr] <= mem_MPORT_472_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_473_en & mem_MPORT_473_mask) begin
      mem[mem_MPORT_473_addr] <= mem_MPORT_473_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_474_en & mem_MPORT_474_mask) begin
      mem[mem_MPORT_474_addr] <= mem_MPORT_474_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_475_en & mem_MPORT_475_mask) begin
      mem[mem_MPORT_475_addr] <= mem_MPORT_475_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_476_en & mem_MPORT_476_mask) begin
      mem[mem_MPORT_476_addr] <= mem_MPORT_476_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_477_en & mem_MPORT_477_mask) begin
      mem[mem_MPORT_477_addr] <= mem_MPORT_477_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_478_en & mem_MPORT_478_mask) begin
      mem[mem_MPORT_478_addr] <= mem_MPORT_478_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_479_en & mem_MPORT_479_mask) begin
      mem[mem_MPORT_479_addr] <= mem_MPORT_479_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_480_en & mem_MPORT_480_mask) begin
      mem[mem_MPORT_480_addr] <= mem_MPORT_480_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_481_en & mem_MPORT_481_mask) begin
      mem[mem_MPORT_481_addr] <= mem_MPORT_481_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_482_en & mem_MPORT_482_mask) begin
      mem[mem_MPORT_482_addr] <= mem_MPORT_482_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_483_en & mem_MPORT_483_mask) begin
      mem[mem_MPORT_483_addr] <= mem_MPORT_483_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_484_en & mem_MPORT_484_mask) begin
      mem[mem_MPORT_484_addr] <= mem_MPORT_484_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_485_en & mem_MPORT_485_mask) begin
      mem[mem_MPORT_485_addr] <= mem_MPORT_485_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_486_en & mem_MPORT_486_mask) begin
      mem[mem_MPORT_486_addr] <= mem_MPORT_486_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_487_en & mem_MPORT_487_mask) begin
      mem[mem_MPORT_487_addr] <= mem_MPORT_487_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_488_en & mem_MPORT_488_mask) begin
      mem[mem_MPORT_488_addr] <= mem_MPORT_488_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_489_en & mem_MPORT_489_mask) begin
      mem[mem_MPORT_489_addr] <= mem_MPORT_489_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_490_en & mem_MPORT_490_mask) begin
      mem[mem_MPORT_490_addr] <= mem_MPORT_490_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_491_en & mem_MPORT_491_mask) begin
      mem[mem_MPORT_491_addr] <= mem_MPORT_491_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_492_en & mem_MPORT_492_mask) begin
      mem[mem_MPORT_492_addr] <= mem_MPORT_492_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_493_en & mem_MPORT_493_mask) begin
      mem[mem_MPORT_493_addr] <= mem_MPORT_493_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_494_en & mem_MPORT_494_mask) begin
      mem[mem_MPORT_494_addr] <= mem_MPORT_494_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_495_en & mem_MPORT_495_mask) begin
      mem[mem_MPORT_495_addr] <= mem_MPORT_495_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_496_en & mem_MPORT_496_mask) begin
      mem[mem_MPORT_496_addr] <= mem_MPORT_496_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_497_en & mem_MPORT_497_mask) begin
      mem[mem_MPORT_497_addr] <= mem_MPORT_497_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_498_en & mem_MPORT_498_mask) begin
      mem[mem_MPORT_498_addr] <= mem_MPORT_498_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_499_en & mem_MPORT_499_mask) begin
      mem[mem_MPORT_499_addr] <= mem_MPORT_499_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_500_en & mem_MPORT_500_mask) begin
      mem[mem_MPORT_500_addr] <= mem_MPORT_500_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_501_en & mem_MPORT_501_mask) begin
      mem[mem_MPORT_501_addr] <= mem_MPORT_501_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_502_en & mem_MPORT_502_mask) begin
      mem[mem_MPORT_502_addr] <= mem_MPORT_502_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_503_en & mem_MPORT_503_mask) begin
      mem[mem_MPORT_503_addr] <= mem_MPORT_503_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_504_en & mem_MPORT_504_mask) begin
      mem[mem_MPORT_504_addr] <= mem_MPORT_504_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_505_en & mem_MPORT_505_mask) begin
      mem[mem_MPORT_505_addr] <= mem_MPORT_505_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_506_en & mem_MPORT_506_mask) begin
      mem[mem_MPORT_506_addr] <= mem_MPORT_506_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_507_en & mem_MPORT_507_mask) begin
      mem[mem_MPORT_507_addr] <= mem_MPORT_507_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_508_en & mem_MPORT_508_mask) begin
      mem[mem_MPORT_508_addr] <= mem_MPORT_508_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_509_en & mem_MPORT_509_mask) begin
      mem[mem_MPORT_509_addr] <= mem_MPORT_509_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_510_en & mem_MPORT_510_mask) begin
      mem[mem_MPORT_510_addr] <= mem_MPORT_510_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_511_en & mem_MPORT_511_mask) begin
      mem[mem_MPORT_511_addr] <= mem_MPORT_511_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_512_en & mem_MPORT_512_mask) begin
      mem[mem_MPORT_512_addr] <= mem_MPORT_512_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem[initvar] = _RAND_0[18:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_14(
  input         clock,
  input         reset,
  input  [8:0]  io_r_addr,
  output [18:0] io_r_data_0,
  output [18:0] io_r_data_1,
  output [18:0] io_r_data_2,
  output [18:0] io_r_data_3,
  input         io_w_en,
  input  [8:0]  io_w_addr,
  input  [18:0] io_w_data_0,
  input  [18:0] io_w_data_1,
  input  [18:0] io_w_data_2,
  input  [18:0] io_w_data_3,
  input  [3:0]  io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [18:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [18:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [18:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [18:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [18:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [18:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [18:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [18:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P_96 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P_96 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P_96 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P_96 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
endmodule
module BankRAM_2P_100(
  input        clock,
  input        reset,
  input  [8:0] io_r_addr,
  output [1:0] io_r_data,
  input        io_w_en,
  input  [8:0] io_w_addr,
  input  [1:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] mem [0:511]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_129_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_130_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_131_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_132_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_133_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_134_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_135_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_136_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_137_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_138_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_139_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_140_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_141_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_142_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_143_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_144_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_145_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_146_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_147_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_148_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_149_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_150_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_151_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_152_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_153_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_154_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_155_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_156_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_157_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_158_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_159_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_160_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_161_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_162_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_163_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_164_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_165_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_166_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_167_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_168_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_169_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_170_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_171_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_172_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_173_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_174_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_175_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_176_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_177_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_178_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_179_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_180_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_181_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_182_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_183_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_184_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_185_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_186_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_187_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_188_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_189_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_190_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_191_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_192_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_193_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_194_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_195_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_196_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_197_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_198_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_199_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_200_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_201_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_202_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_203_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_204_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_205_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_206_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_207_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_208_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_209_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_210_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_211_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_212_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_213_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_214_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_215_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_216_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_217_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_218_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_219_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_220_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_221_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_222_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_223_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_224_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_225_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_226_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_227_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_228_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_229_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_230_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_231_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_232_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_233_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_234_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_235_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_236_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_237_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_238_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_239_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_240_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_241_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_242_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_243_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_244_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_245_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_246_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_247_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_248_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_249_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_250_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_251_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_252_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_253_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_254_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_255_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_256_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_257_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_257_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_257_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_257_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_258_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_258_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_258_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_258_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_259_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_259_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_259_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_259_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_260_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_260_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_260_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_260_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_261_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_261_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_261_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_261_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_262_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_262_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_262_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_262_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_263_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_263_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_263_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_263_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_264_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_264_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_264_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_264_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_265_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_265_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_265_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_265_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_266_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_266_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_266_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_266_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_267_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_267_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_267_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_267_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_268_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_268_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_268_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_268_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_269_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_269_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_269_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_269_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_270_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_270_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_270_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_270_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_271_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_271_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_271_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_271_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_272_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_272_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_272_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_272_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_273_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_273_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_273_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_273_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_274_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_274_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_274_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_274_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_275_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_275_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_275_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_275_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_276_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_276_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_276_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_276_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_277_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_277_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_277_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_277_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_278_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_278_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_278_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_278_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_279_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_279_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_279_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_279_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_280_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_280_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_280_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_280_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_281_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_281_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_281_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_281_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_282_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_282_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_282_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_282_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_283_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_283_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_283_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_283_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_284_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_284_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_284_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_284_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_285_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_285_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_285_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_285_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_286_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_286_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_286_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_286_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_287_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_287_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_287_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_287_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_288_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_288_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_288_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_288_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_289_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_289_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_289_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_289_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_290_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_290_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_290_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_290_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_291_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_291_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_291_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_291_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_292_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_292_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_292_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_292_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_293_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_293_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_293_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_293_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_294_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_294_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_294_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_294_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_295_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_295_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_295_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_295_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_296_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_296_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_296_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_296_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_297_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_297_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_297_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_297_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_298_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_298_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_298_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_298_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_299_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_299_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_299_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_299_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_300_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_300_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_300_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_300_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_301_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_301_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_301_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_301_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_302_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_302_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_302_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_302_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_303_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_303_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_303_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_303_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_304_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_304_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_304_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_304_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_305_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_305_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_305_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_305_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_306_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_306_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_306_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_306_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_307_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_307_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_307_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_307_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_308_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_308_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_308_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_308_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_309_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_309_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_309_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_309_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_310_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_310_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_310_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_310_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_311_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_311_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_311_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_311_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_312_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_312_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_312_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_312_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_313_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_313_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_313_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_313_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_314_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_314_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_314_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_314_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_315_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_315_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_315_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_315_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_316_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_316_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_316_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_316_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_317_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_317_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_317_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_317_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_318_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_318_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_318_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_318_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_319_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_319_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_319_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_319_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_320_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_320_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_320_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_320_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_321_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_321_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_321_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_321_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_322_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_322_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_322_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_322_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_323_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_323_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_323_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_323_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_324_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_324_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_324_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_324_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_325_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_325_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_325_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_325_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_326_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_326_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_326_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_326_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_327_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_327_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_327_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_327_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_328_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_328_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_328_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_328_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_329_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_329_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_329_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_329_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_330_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_330_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_330_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_330_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_331_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_331_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_331_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_331_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_332_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_332_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_332_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_332_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_333_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_333_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_333_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_333_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_334_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_334_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_334_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_334_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_335_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_335_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_335_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_335_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_336_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_336_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_336_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_336_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_337_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_337_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_337_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_337_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_338_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_338_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_338_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_338_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_339_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_339_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_339_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_339_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_340_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_340_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_340_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_340_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_341_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_341_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_341_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_341_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_342_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_342_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_342_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_342_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_343_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_343_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_343_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_343_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_344_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_344_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_344_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_344_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_345_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_345_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_345_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_345_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_346_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_346_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_346_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_346_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_347_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_347_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_347_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_347_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_348_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_348_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_348_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_348_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_349_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_349_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_349_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_349_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_350_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_350_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_350_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_350_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_351_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_351_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_351_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_351_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_352_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_352_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_352_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_352_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_353_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_353_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_353_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_353_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_354_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_354_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_354_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_354_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_355_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_355_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_355_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_355_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_356_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_356_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_356_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_356_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_357_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_357_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_357_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_357_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_358_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_358_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_358_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_358_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_359_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_359_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_359_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_359_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_360_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_360_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_360_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_360_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_361_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_361_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_361_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_361_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_362_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_362_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_362_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_362_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_363_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_363_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_363_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_363_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_364_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_364_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_364_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_364_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_365_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_365_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_365_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_365_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_366_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_366_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_366_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_366_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_367_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_367_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_367_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_367_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_368_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_368_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_368_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_368_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_369_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_369_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_369_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_369_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_370_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_370_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_370_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_370_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_371_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_371_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_371_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_371_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_372_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_372_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_372_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_372_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_373_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_373_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_373_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_373_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_374_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_374_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_374_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_374_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_375_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_375_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_375_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_375_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_376_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_376_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_376_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_376_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_377_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_377_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_377_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_377_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_378_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_378_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_378_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_378_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_379_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_379_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_379_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_379_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_380_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_380_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_380_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_380_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_381_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_381_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_381_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_381_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_382_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_382_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_382_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_382_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_383_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_383_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_383_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_383_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_384_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_384_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_384_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_384_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_385_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_385_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_385_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_385_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_386_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_386_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_386_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_386_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_387_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_387_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_387_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_387_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_388_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_388_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_388_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_388_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_389_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_389_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_389_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_389_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_390_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_390_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_390_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_390_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_391_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_391_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_391_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_391_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_392_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_392_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_392_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_392_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_393_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_393_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_393_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_393_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_394_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_394_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_394_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_394_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_395_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_395_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_395_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_395_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_396_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_396_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_396_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_396_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_397_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_397_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_397_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_397_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_398_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_398_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_398_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_398_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_399_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_399_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_399_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_399_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_400_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_400_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_400_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_400_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_401_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_401_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_401_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_401_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_402_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_402_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_402_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_402_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_403_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_403_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_403_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_403_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_404_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_404_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_404_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_404_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_405_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_405_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_405_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_405_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_406_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_406_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_406_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_406_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_407_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_407_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_407_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_407_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_408_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_408_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_408_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_408_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_409_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_409_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_409_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_409_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_410_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_410_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_410_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_410_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_411_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_411_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_411_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_411_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_412_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_412_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_412_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_412_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_413_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_413_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_413_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_413_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_414_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_414_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_414_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_414_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_415_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_415_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_415_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_415_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_416_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_416_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_416_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_416_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_417_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_417_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_417_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_417_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_418_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_418_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_418_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_418_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_419_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_419_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_419_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_419_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_420_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_420_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_420_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_420_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_421_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_421_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_421_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_421_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_422_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_422_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_422_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_422_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_423_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_423_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_423_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_423_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_424_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_424_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_424_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_424_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_425_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_425_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_425_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_425_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_426_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_426_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_426_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_426_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_427_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_427_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_427_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_427_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_428_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_428_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_428_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_428_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_429_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_429_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_429_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_429_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_430_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_430_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_430_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_430_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_431_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_431_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_431_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_431_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_432_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_432_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_432_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_432_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_433_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_433_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_433_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_433_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_434_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_434_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_434_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_434_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_435_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_435_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_435_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_435_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_436_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_436_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_436_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_436_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_437_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_437_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_437_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_437_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_438_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_438_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_438_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_438_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_439_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_439_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_439_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_439_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_440_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_440_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_440_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_440_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_441_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_441_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_441_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_441_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_442_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_442_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_442_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_442_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_443_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_443_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_443_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_443_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_444_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_444_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_444_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_444_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_445_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_445_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_445_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_445_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_446_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_446_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_446_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_446_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_447_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_447_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_447_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_447_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_448_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_448_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_448_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_448_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_449_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_449_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_449_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_449_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_450_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_450_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_450_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_450_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_451_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_451_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_451_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_451_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_452_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_452_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_452_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_452_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_453_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_453_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_453_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_453_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_454_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_454_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_454_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_454_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_455_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_455_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_455_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_455_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_456_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_456_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_456_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_456_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_457_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_457_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_457_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_457_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_458_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_458_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_458_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_458_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_459_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_459_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_459_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_459_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_460_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_460_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_460_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_460_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_461_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_461_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_461_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_461_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_462_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_462_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_462_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_462_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_463_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_463_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_463_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_463_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_464_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_464_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_464_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_464_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_465_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_465_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_465_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_465_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_466_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_466_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_466_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_466_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_467_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_467_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_467_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_467_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_468_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_468_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_468_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_468_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_469_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_469_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_469_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_469_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_470_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_470_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_470_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_470_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_471_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_471_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_471_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_471_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_472_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_472_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_472_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_472_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_473_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_473_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_473_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_473_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_474_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_474_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_474_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_474_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_475_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_475_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_475_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_475_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_476_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_476_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_476_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_476_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_477_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_477_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_477_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_477_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_478_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_478_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_478_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_478_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_479_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_479_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_479_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_479_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_480_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_480_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_480_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_480_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_481_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_481_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_481_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_481_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_482_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_482_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_482_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_482_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_483_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_483_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_483_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_483_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_484_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_484_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_484_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_484_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_485_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_485_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_485_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_485_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_486_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_486_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_486_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_486_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_487_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_487_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_487_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_487_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_488_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_488_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_488_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_488_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_489_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_489_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_489_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_489_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_490_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_490_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_490_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_490_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_491_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_491_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_491_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_491_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_492_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_492_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_492_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_492_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_493_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_493_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_493_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_493_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_494_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_494_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_494_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_494_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_495_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_495_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_495_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_495_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_496_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_496_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_496_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_496_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_497_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_497_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_497_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_497_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_498_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_498_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_498_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_498_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_499_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_499_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_499_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_499_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_500_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_500_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_500_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_500_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_501_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_501_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_501_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_501_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_502_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_502_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_502_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_502_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_503_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_503_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_503_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_503_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_504_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_504_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_504_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_504_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_505_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_505_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_505_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_505_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_506_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_506_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_506_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_506_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_507_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_507_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_507_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_507_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_508_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_508_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_508_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_508_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_509_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_509_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_509_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_509_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_510_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_510_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_510_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_510_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_511_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_511_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_511_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_511_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_512_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_512_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_512_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_512_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [8:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 2'h0;
  assign mem_MPORT_addr = 9'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 2'h0;
  assign mem_MPORT_1_addr = 9'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 2'h0;
  assign mem_MPORT_2_addr = 9'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 2'h0;
  assign mem_MPORT_3_addr = 9'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 2'h0;
  assign mem_MPORT_4_addr = 9'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 2'h0;
  assign mem_MPORT_5_addr = 9'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 2'h0;
  assign mem_MPORT_6_addr = 9'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 2'h0;
  assign mem_MPORT_7_addr = 9'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 2'h0;
  assign mem_MPORT_8_addr = 9'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 2'h0;
  assign mem_MPORT_9_addr = 9'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 2'h0;
  assign mem_MPORT_10_addr = 9'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 2'h0;
  assign mem_MPORT_11_addr = 9'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 2'h0;
  assign mem_MPORT_12_addr = 9'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 2'h0;
  assign mem_MPORT_13_addr = 9'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 2'h0;
  assign mem_MPORT_14_addr = 9'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 2'h0;
  assign mem_MPORT_15_addr = 9'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 2'h0;
  assign mem_MPORT_16_addr = 9'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 2'h0;
  assign mem_MPORT_17_addr = 9'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 2'h0;
  assign mem_MPORT_18_addr = 9'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 2'h0;
  assign mem_MPORT_19_addr = 9'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 2'h0;
  assign mem_MPORT_20_addr = 9'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 2'h0;
  assign mem_MPORT_21_addr = 9'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 2'h0;
  assign mem_MPORT_22_addr = 9'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 2'h0;
  assign mem_MPORT_23_addr = 9'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 2'h0;
  assign mem_MPORT_24_addr = 9'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 2'h0;
  assign mem_MPORT_25_addr = 9'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 2'h0;
  assign mem_MPORT_26_addr = 9'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 2'h0;
  assign mem_MPORT_27_addr = 9'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 2'h0;
  assign mem_MPORT_28_addr = 9'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 2'h0;
  assign mem_MPORT_29_addr = 9'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 2'h0;
  assign mem_MPORT_30_addr = 9'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 2'h0;
  assign mem_MPORT_31_addr = 9'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 2'h0;
  assign mem_MPORT_32_addr = 9'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 2'h0;
  assign mem_MPORT_33_addr = 9'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 2'h0;
  assign mem_MPORT_34_addr = 9'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 2'h0;
  assign mem_MPORT_35_addr = 9'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 2'h0;
  assign mem_MPORT_36_addr = 9'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 2'h0;
  assign mem_MPORT_37_addr = 9'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 2'h0;
  assign mem_MPORT_38_addr = 9'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 2'h0;
  assign mem_MPORT_39_addr = 9'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 2'h0;
  assign mem_MPORT_40_addr = 9'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 2'h0;
  assign mem_MPORT_41_addr = 9'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 2'h0;
  assign mem_MPORT_42_addr = 9'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 2'h0;
  assign mem_MPORT_43_addr = 9'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 2'h0;
  assign mem_MPORT_44_addr = 9'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 2'h0;
  assign mem_MPORT_45_addr = 9'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 2'h0;
  assign mem_MPORT_46_addr = 9'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 2'h0;
  assign mem_MPORT_47_addr = 9'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 2'h0;
  assign mem_MPORT_48_addr = 9'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 2'h0;
  assign mem_MPORT_49_addr = 9'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 2'h0;
  assign mem_MPORT_50_addr = 9'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 2'h0;
  assign mem_MPORT_51_addr = 9'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 2'h0;
  assign mem_MPORT_52_addr = 9'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 2'h0;
  assign mem_MPORT_53_addr = 9'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 2'h0;
  assign mem_MPORT_54_addr = 9'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 2'h0;
  assign mem_MPORT_55_addr = 9'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 2'h0;
  assign mem_MPORT_56_addr = 9'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 2'h0;
  assign mem_MPORT_57_addr = 9'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 2'h0;
  assign mem_MPORT_58_addr = 9'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 2'h0;
  assign mem_MPORT_59_addr = 9'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 2'h0;
  assign mem_MPORT_60_addr = 9'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 2'h0;
  assign mem_MPORT_61_addr = 9'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 2'h0;
  assign mem_MPORT_62_addr = 9'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 2'h0;
  assign mem_MPORT_63_addr = 9'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 2'h0;
  assign mem_MPORT_64_addr = 9'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 2'h0;
  assign mem_MPORT_65_addr = 9'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 2'h0;
  assign mem_MPORT_66_addr = 9'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 2'h0;
  assign mem_MPORT_67_addr = 9'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 2'h0;
  assign mem_MPORT_68_addr = 9'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 2'h0;
  assign mem_MPORT_69_addr = 9'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 2'h0;
  assign mem_MPORT_70_addr = 9'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 2'h0;
  assign mem_MPORT_71_addr = 9'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 2'h0;
  assign mem_MPORT_72_addr = 9'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 2'h0;
  assign mem_MPORT_73_addr = 9'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 2'h0;
  assign mem_MPORT_74_addr = 9'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 2'h0;
  assign mem_MPORT_75_addr = 9'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 2'h0;
  assign mem_MPORT_76_addr = 9'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 2'h0;
  assign mem_MPORT_77_addr = 9'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 2'h0;
  assign mem_MPORT_78_addr = 9'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 2'h0;
  assign mem_MPORT_79_addr = 9'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 2'h0;
  assign mem_MPORT_80_addr = 9'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 2'h0;
  assign mem_MPORT_81_addr = 9'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 2'h0;
  assign mem_MPORT_82_addr = 9'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 2'h0;
  assign mem_MPORT_83_addr = 9'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 2'h0;
  assign mem_MPORT_84_addr = 9'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 2'h0;
  assign mem_MPORT_85_addr = 9'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 2'h0;
  assign mem_MPORT_86_addr = 9'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 2'h0;
  assign mem_MPORT_87_addr = 9'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 2'h0;
  assign mem_MPORT_88_addr = 9'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 2'h0;
  assign mem_MPORT_89_addr = 9'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 2'h0;
  assign mem_MPORT_90_addr = 9'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 2'h0;
  assign mem_MPORT_91_addr = 9'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 2'h0;
  assign mem_MPORT_92_addr = 9'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 2'h0;
  assign mem_MPORT_93_addr = 9'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 2'h0;
  assign mem_MPORT_94_addr = 9'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 2'h0;
  assign mem_MPORT_95_addr = 9'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 2'h0;
  assign mem_MPORT_96_addr = 9'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 2'h0;
  assign mem_MPORT_97_addr = 9'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 2'h0;
  assign mem_MPORT_98_addr = 9'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 2'h0;
  assign mem_MPORT_99_addr = 9'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 2'h0;
  assign mem_MPORT_100_addr = 9'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 2'h0;
  assign mem_MPORT_101_addr = 9'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 2'h0;
  assign mem_MPORT_102_addr = 9'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 2'h0;
  assign mem_MPORT_103_addr = 9'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 2'h0;
  assign mem_MPORT_104_addr = 9'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 2'h0;
  assign mem_MPORT_105_addr = 9'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 2'h0;
  assign mem_MPORT_106_addr = 9'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 2'h0;
  assign mem_MPORT_107_addr = 9'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 2'h0;
  assign mem_MPORT_108_addr = 9'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 2'h0;
  assign mem_MPORT_109_addr = 9'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 2'h0;
  assign mem_MPORT_110_addr = 9'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 2'h0;
  assign mem_MPORT_111_addr = 9'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 2'h0;
  assign mem_MPORT_112_addr = 9'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 2'h0;
  assign mem_MPORT_113_addr = 9'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 2'h0;
  assign mem_MPORT_114_addr = 9'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 2'h0;
  assign mem_MPORT_115_addr = 9'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 2'h0;
  assign mem_MPORT_116_addr = 9'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 2'h0;
  assign mem_MPORT_117_addr = 9'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 2'h0;
  assign mem_MPORT_118_addr = 9'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 2'h0;
  assign mem_MPORT_119_addr = 9'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 2'h0;
  assign mem_MPORT_120_addr = 9'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 2'h0;
  assign mem_MPORT_121_addr = 9'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 2'h0;
  assign mem_MPORT_122_addr = 9'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 2'h0;
  assign mem_MPORT_123_addr = 9'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 2'h0;
  assign mem_MPORT_124_addr = 9'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 2'h0;
  assign mem_MPORT_125_addr = 9'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 2'h0;
  assign mem_MPORT_126_addr = 9'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 2'h0;
  assign mem_MPORT_127_addr = 9'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 2'h0;
  assign mem_MPORT_128_addr = 9'h80;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = reset;
  assign mem_MPORT_129_data = 2'h0;
  assign mem_MPORT_129_addr = 9'h81;
  assign mem_MPORT_129_mask = 1'h1;
  assign mem_MPORT_129_en = reset;
  assign mem_MPORT_130_data = 2'h0;
  assign mem_MPORT_130_addr = 9'h82;
  assign mem_MPORT_130_mask = 1'h1;
  assign mem_MPORT_130_en = reset;
  assign mem_MPORT_131_data = 2'h0;
  assign mem_MPORT_131_addr = 9'h83;
  assign mem_MPORT_131_mask = 1'h1;
  assign mem_MPORT_131_en = reset;
  assign mem_MPORT_132_data = 2'h0;
  assign mem_MPORT_132_addr = 9'h84;
  assign mem_MPORT_132_mask = 1'h1;
  assign mem_MPORT_132_en = reset;
  assign mem_MPORT_133_data = 2'h0;
  assign mem_MPORT_133_addr = 9'h85;
  assign mem_MPORT_133_mask = 1'h1;
  assign mem_MPORT_133_en = reset;
  assign mem_MPORT_134_data = 2'h0;
  assign mem_MPORT_134_addr = 9'h86;
  assign mem_MPORT_134_mask = 1'h1;
  assign mem_MPORT_134_en = reset;
  assign mem_MPORT_135_data = 2'h0;
  assign mem_MPORT_135_addr = 9'h87;
  assign mem_MPORT_135_mask = 1'h1;
  assign mem_MPORT_135_en = reset;
  assign mem_MPORT_136_data = 2'h0;
  assign mem_MPORT_136_addr = 9'h88;
  assign mem_MPORT_136_mask = 1'h1;
  assign mem_MPORT_136_en = reset;
  assign mem_MPORT_137_data = 2'h0;
  assign mem_MPORT_137_addr = 9'h89;
  assign mem_MPORT_137_mask = 1'h1;
  assign mem_MPORT_137_en = reset;
  assign mem_MPORT_138_data = 2'h0;
  assign mem_MPORT_138_addr = 9'h8a;
  assign mem_MPORT_138_mask = 1'h1;
  assign mem_MPORT_138_en = reset;
  assign mem_MPORT_139_data = 2'h0;
  assign mem_MPORT_139_addr = 9'h8b;
  assign mem_MPORT_139_mask = 1'h1;
  assign mem_MPORT_139_en = reset;
  assign mem_MPORT_140_data = 2'h0;
  assign mem_MPORT_140_addr = 9'h8c;
  assign mem_MPORT_140_mask = 1'h1;
  assign mem_MPORT_140_en = reset;
  assign mem_MPORT_141_data = 2'h0;
  assign mem_MPORT_141_addr = 9'h8d;
  assign mem_MPORT_141_mask = 1'h1;
  assign mem_MPORT_141_en = reset;
  assign mem_MPORT_142_data = 2'h0;
  assign mem_MPORT_142_addr = 9'h8e;
  assign mem_MPORT_142_mask = 1'h1;
  assign mem_MPORT_142_en = reset;
  assign mem_MPORT_143_data = 2'h0;
  assign mem_MPORT_143_addr = 9'h8f;
  assign mem_MPORT_143_mask = 1'h1;
  assign mem_MPORT_143_en = reset;
  assign mem_MPORT_144_data = 2'h0;
  assign mem_MPORT_144_addr = 9'h90;
  assign mem_MPORT_144_mask = 1'h1;
  assign mem_MPORT_144_en = reset;
  assign mem_MPORT_145_data = 2'h0;
  assign mem_MPORT_145_addr = 9'h91;
  assign mem_MPORT_145_mask = 1'h1;
  assign mem_MPORT_145_en = reset;
  assign mem_MPORT_146_data = 2'h0;
  assign mem_MPORT_146_addr = 9'h92;
  assign mem_MPORT_146_mask = 1'h1;
  assign mem_MPORT_146_en = reset;
  assign mem_MPORT_147_data = 2'h0;
  assign mem_MPORT_147_addr = 9'h93;
  assign mem_MPORT_147_mask = 1'h1;
  assign mem_MPORT_147_en = reset;
  assign mem_MPORT_148_data = 2'h0;
  assign mem_MPORT_148_addr = 9'h94;
  assign mem_MPORT_148_mask = 1'h1;
  assign mem_MPORT_148_en = reset;
  assign mem_MPORT_149_data = 2'h0;
  assign mem_MPORT_149_addr = 9'h95;
  assign mem_MPORT_149_mask = 1'h1;
  assign mem_MPORT_149_en = reset;
  assign mem_MPORT_150_data = 2'h0;
  assign mem_MPORT_150_addr = 9'h96;
  assign mem_MPORT_150_mask = 1'h1;
  assign mem_MPORT_150_en = reset;
  assign mem_MPORT_151_data = 2'h0;
  assign mem_MPORT_151_addr = 9'h97;
  assign mem_MPORT_151_mask = 1'h1;
  assign mem_MPORT_151_en = reset;
  assign mem_MPORT_152_data = 2'h0;
  assign mem_MPORT_152_addr = 9'h98;
  assign mem_MPORT_152_mask = 1'h1;
  assign mem_MPORT_152_en = reset;
  assign mem_MPORT_153_data = 2'h0;
  assign mem_MPORT_153_addr = 9'h99;
  assign mem_MPORT_153_mask = 1'h1;
  assign mem_MPORT_153_en = reset;
  assign mem_MPORT_154_data = 2'h0;
  assign mem_MPORT_154_addr = 9'h9a;
  assign mem_MPORT_154_mask = 1'h1;
  assign mem_MPORT_154_en = reset;
  assign mem_MPORT_155_data = 2'h0;
  assign mem_MPORT_155_addr = 9'h9b;
  assign mem_MPORT_155_mask = 1'h1;
  assign mem_MPORT_155_en = reset;
  assign mem_MPORT_156_data = 2'h0;
  assign mem_MPORT_156_addr = 9'h9c;
  assign mem_MPORT_156_mask = 1'h1;
  assign mem_MPORT_156_en = reset;
  assign mem_MPORT_157_data = 2'h0;
  assign mem_MPORT_157_addr = 9'h9d;
  assign mem_MPORT_157_mask = 1'h1;
  assign mem_MPORT_157_en = reset;
  assign mem_MPORT_158_data = 2'h0;
  assign mem_MPORT_158_addr = 9'h9e;
  assign mem_MPORT_158_mask = 1'h1;
  assign mem_MPORT_158_en = reset;
  assign mem_MPORT_159_data = 2'h0;
  assign mem_MPORT_159_addr = 9'h9f;
  assign mem_MPORT_159_mask = 1'h1;
  assign mem_MPORT_159_en = reset;
  assign mem_MPORT_160_data = 2'h0;
  assign mem_MPORT_160_addr = 9'ha0;
  assign mem_MPORT_160_mask = 1'h1;
  assign mem_MPORT_160_en = reset;
  assign mem_MPORT_161_data = 2'h0;
  assign mem_MPORT_161_addr = 9'ha1;
  assign mem_MPORT_161_mask = 1'h1;
  assign mem_MPORT_161_en = reset;
  assign mem_MPORT_162_data = 2'h0;
  assign mem_MPORT_162_addr = 9'ha2;
  assign mem_MPORT_162_mask = 1'h1;
  assign mem_MPORT_162_en = reset;
  assign mem_MPORT_163_data = 2'h0;
  assign mem_MPORT_163_addr = 9'ha3;
  assign mem_MPORT_163_mask = 1'h1;
  assign mem_MPORT_163_en = reset;
  assign mem_MPORT_164_data = 2'h0;
  assign mem_MPORT_164_addr = 9'ha4;
  assign mem_MPORT_164_mask = 1'h1;
  assign mem_MPORT_164_en = reset;
  assign mem_MPORT_165_data = 2'h0;
  assign mem_MPORT_165_addr = 9'ha5;
  assign mem_MPORT_165_mask = 1'h1;
  assign mem_MPORT_165_en = reset;
  assign mem_MPORT_166_data = 2'h0;
  assign mem_MPORT_166_addr = 9'ha6;
  assign mem_MPORT_166_mask = 1'h1;
  assign mem_MPORT_166_en = reset;
  assign mem_MPORT_167_data = 2'h0;
  assign mem_MPORT_167_addr = 9'ha7;
  assign mem_MPORT_167_mask = 1'h1;
  assign mem_MPORT_167_en = reset;
  assign mem_MPORT_168_data = 2'h0;
  assign mem_MPORT_168_addr = 9'ha8;
  assign mem_MPORT_168_mask = 1'h1;
  assign mem_MPORT_168_en = reset;
  assign mem_MPORT_169_data = 2'h0;
  assign mem_MPORT_169_addr = 9'ha9;
  assign mem_MPORT_169_mask = 1'h1;
  assign mem_MPORT_169_en = reset;
  assign mem_MPORT_170_data = 2'h0;
  assign mem_MPORT_170_addr = 9'haa;
  assign mem_MPORT_170_mask = 1'h1;
  assign mem_MPORT_170_en = reset;
  assign mem_MPORT_171_data = 2'h0;
  assign mem_MPORT_171_addr = 9'hab;
  assign mem_MPORT_171_mask = 1'h1;
  assign mem_MPORT_171_en = reset;
  assign mem_MPORT_172_data = 2'h0;
  assign mem_MPORT_172_addr = 9'hac;
  assign mem_MPORT_172_mask = 1'h1;
  assign mem_MPORT_172_en = reset;
  assign mem_MPORT_173_data = 2'h0;
  assign mem_MPORT_173_addr = 9'had;
  assign mem_MPORT_173_mask = 1'h1;
  assign mem_MPORT_173_en = reset;
  assign mem_MPORT_174_data = 2'h0;
  assign mem_MPORT_174_addr = 9'hae;
  assign mem_MPORT_174_mask = 1'h1;
  assign mem_MPORT_174_en = reset;
  assign mem_MPORT_175_data = 2'h0;
  assign mem_MPORT_175_addr = 9'haf;
  assign mem_MPORT_175_mask = 1'h1;
  assign mem_MPORT_175_en = reset;
  assign mem_MPORT_176_data = 2'h0;
  assign mem_MPORT_176_addr = 9'hb0;
  assign mem_MPORT_176_mask = 1'h1;
  assign mem_MPORT_176_en = reset;
  assign mem_MPORT_177_data = 2'h0;
  assign mem_MPORT_177_addr = 9'hb1;
  assign mem_MPORT_177_mask = 1'h1;
  assign mem_MPORT_177_en = reset;
  assign mem_MPORT_178_data = 2'h0;
  assign mem_MPORT_178_addr = 9'hb2;
  assign mem_MPORT_178_mask = 1'h1;
  assign mem_MPORT_178_en = reset;
  assign mem_MPORT_179_data = 2'h0;
  assign mem_MPORT_179_addr = 9'hb3;
  assign mem_MPORT_179_mask = 1'h1;
  assign mem_MPORT_179_en = reset;
  assign mem_MPORT_180_data = 2'h0;
  assign mem_MPORT_180_addr = 9'hb4;
  assign mem_MPORT_180_mask = 1'h1;
  assign mem_MPORT_180_en = reset;
  assign mem_MPORT_181_data = 2'h0;
  assign mem_MPORT_181_addr = 9'hb5;
  assign mem_MPORT_181_mask = 1'h1;
  assign mem_MPORT_181_en = reset;
  assign mem_MPORT_182_data = 2'h0;
  assign mem_MPORT_182_addr = 9'hb6;
  assign mem_MPORT_182_mask = 1'h1;
  assign mem_MPORT_182_en = reset;
  assign mem_MPORT_183_data = 2'h0;
  assign mem_MPORT_183_addr = 9'hb7;
  assign mem_MPORT_183_mask = 1'h1;
  assign mem_MPORT_183_en = reset;
  assign mem_MPORT_184_data = 2'h0;
  assign mem_MPORT_184_addr = 9'hb8;
  assign mem_MPORT_184_mask = 1'h1;
  assign mem_MPORT_184_en = reset;
  assign mem_MPORT_185_data = 2'h0;
  assign mem_MPORT_185_addr = 9'hb9;
  assign mem_MPORT_185_mask = 1'h1;
  assign mem_MPORT_185_en = reset;
  assign mem_MPORT_186_data = 2'h0;
  assign mem_MPORT_186_addr = 9'hba;
  assign mem_MPORT_186_mask = 1'h1;
  assign mem_MPORT_186_en = reset;
  assign mem_MPORT_187_data = 2'h0;
  assign mem_MPORT_187_addr = 9'hbb;
  assign mem_MPORT_187_mask = 1'h1;
  assign mem_MPORT_187_en = reset;
  assign mem_MPORT_188_data = 2'h0;
  assign mem_MPORT_188_addr = 9'hbc;
  assign mem_MPORT_188_mask = 1'h1;
  assign mem_MPORT_188_en = reset;
  assign mem_MPORT_189_data = 2'h0;
  assign mem_MPORT_189_addr = 9'hbd;
  assign mem_MPORT_189_mask = 1'h1;
  assign mem_MPORT_189_en = reset;
  assign mem_MPORT_190_data = 2'h0;
  assign mem_MPORT_190_addr = 9'hbe;
  assign mem_MPORT_190_mask = 1'h1;
  assign mem_MPORT_190_en = reset;
  assign mem_MPORT_191_data = 2'h0;
  assign mem_MPORT_191_addr = 9'hbf;
  assign mem_MPORT_191_mask = 1'h1;
  assign mem_MPORT_191_en = reset;
  assign mem_MPORT_192_data = 2'h0;
  assign mem_MPORT_192_addr = 9'hc0;
  assign mem_MPORT_192_mask = 1'h1;
  assign mem_MPORT_192_en = reset;
  assign mem_MPORT_193_data = 2'h0;
  assign mem_MPORT_193_addr = 9'hc1;
  assign mem_MPORT_193_mask = 1'h1;
  assign mem_MPORT_193_en = reset;
  assign mem_MPORT_194_data = 2'h0;
  assign mem_MPORT_194_addr = 9'hc2;
  assign mem_MPORT_194_mask = 1'h1;
  assign mem_MPORT_194_en = reset;
  assign mem_MPORT_195_data = 2'h0;
  assign mem_MPORT_195_addr = 9'hc3;
  assign mem_MPORT_195_mask = 1'h1;
  assign mem_MPORT_195_en = reset;
  assign mem_MPORT_196_data = 2'h0;
  assign mem_MPORT_196_addr = 9'hc4;
  assign mem_MPORT_196_mask = 1'h1;
  assign mem_MPORT_196_en = reset;
  assign mem_MPORT_197_data = 2'h0;
  assign mem_MPORT_197_addr = 9'hc5;
  assign mem_MPORT_197_mask = 1'h1;
  assign mem_MPORT_197_en = reset;
  assign mem_MPORT_198_data = 2'h0;
  assign mem_MPORT_198_addr = 9'hc6;
  assign mem_MPORT_198_mask = 1'h1;
  assign mem_MPORT_198_en = reset;
  assign mem_MPORT_199_data = 2'h0;
  assign mem_MPORT_199_addr = 9'hc7;
  assign mem_MPORT_199_mask = 1'h1;
  assign mem_MPORT_199_en = reset;
  assign mem_MPORT_200_data = 2'h0;
  assign mem_MPORT_200_addr = 9'hc8;
  assign mem_MPORT_200_mask = 1'h1;
  assign mem_MPORT_200_en = reset;
  assign mem_MPORT_201_data = 2'h0;
  assign mem_MPORT_201_addr = 9'hc9;
  assign mem_MPORT_201_mask = 1'h1;
  assign mem_MPORT_201_en = reset;
  assign mem_MPORT_202_data = 2'h0;
  assign mem_MPORT_202_addr = 9'hca;
  assign mem_MPORT_202_mask = 1'h1;
  assign mem_MPORT_202_en = reset;
  assign mem_MPORT_203_data = 2'h0;
  assign mem_MPORT_203_addr = 9'hcb;
  assign mem_MPORT_203_mask = 1'h1;
  assign mem_MPORT_203_en = reset;
  assign mem_MPORT_204_data = 2'h0;
  assign mem_MPORT_204_addr = 9'hcc;
  assign mem_MPORT_204_mask = 1'h1;
  assign mem_MPORT_204_en = reset;
  assign mem_MPORT_205_data = 2'h0;
  assign mem_MPORT_205_addr = 9'hcd;
  assign mem_MPORT_205_mask = 1'h1;
  assign mem_MPORT_205_en = reset;
  assign mem_MPORT_206_data = 2'h0;
  assign mem_MPORT_206_addr = 9'hce;
  assign mem_MPORT_206_mask = 1'h1;
  assign mem_MPORT_206_en = reset;
  assign mem_MPORT_207_data = 2'h0;
  assign mem_MPORT_207_addr = 9'hcf;
  assign mem_MPORT_207_mask = 1'h1;
  assign mem_MPORT_207_en = reset;
  assign mem_MPORT_208_data = 2'h0;
  assign mem_MPORT_208_addr = 9'hd0;
  assign mem_MPORT_208_mask = 1'h1;
  assign mem_MPORT_208_en = reset;
  assign mem_MPORT_209_data = 2'h0;
  assign mem_MPORT_209_addr = 9'hd1;
  assign mem_MPORT_209_mask = 1'h1;
  assign mem_MPORT_209_en = reset;
  assign mem_MPORT_210_data = 2'h0;
  assign mem_MPORT_210_addr = 9'hd2;
  assign mem_MPORT_210_mask = 1'h1;
  assign mem_MPORT_210_en = reset;
  assign mem_MPORT_211_data = 2'h0;
  assign mem_MPORT_211_addr = 9'hd3;
  assign mem_MPORT_211_mask = 1'h1;
  assign mem_MPORT_211_en = reset;
  assign mem_MPORT_212_data = 2'h0;
  assign mem_MPORT_212_addr = 9'hd4;
  assign mem_MPORT_212_mask = 1'h1;
  assign mem_MPORT_212_en = reset;
  assign mem_MPORT_213_data = 2'h0;
  assign mem_MPORT_213_addr = 9'hd5;
  assign mem_MPORT_213_mask = 1'h1;
  assign mem_MPORT_213_en = reset;
  assign mem_MPORT_214_data = 2'h0;
  assign mem_MPORT_214_addr = 9'hd6;
  assign mem_MPORT_214_mask = 1'h1;
  assign mem_MPORT_214_en = reset;
  assign mem_MPORT_215_data = 2'h0;
  assign mem_MPORT_215_addr = 9'hd7;
  assign mem_MPORT_215_mask = 1'h1;
  assign mem_MPORT_215_en = reset;
  assign mem_MPORT_216_data = 2'h0;
  assign mem_MPORT_216_addr = 9'hd8;
  assign mem_MPORT_216_mask = 1'h1;
  assign mem_MPORT_216_en = reset;
  assign mem_MPORT_217_data = 2'h0;
  assign mem_MPORT_217_addr = 9'hd9;
  assign mem_MPORT_217_mask = 1'h1;
  assign mem_MPORT_217_en = reset;
  assign mem_MPORT_218_data = 2'h0;
  assign mem_MPORT_218_addr = 9'hda;
  assign mem_MPORT_218_mask = 1'h1;
  assign mem_MPORT_218_en = reset;
  assign mem_MPORT_219_data = 2'h0;
  assign mem_MPORT_219_addr = 9'hdb;
  assign mem_MPORT_219_mask = 1'h1;
  assign mem_MPORT_219_en = reset;
  assign mem_MPORT_220_data = 2'h0;
  assign mem_MPORT_220_addr = 9'hdc;
  assign mem_MPORT_220_mask = 1'h1;
  assign mem_MPORT_220_en = reset;
  assign mem_MPORT_221_data = 2'h0;
  assign mem_MPORT_221_addr = 9'hdd;
  assign mem_MPORT_221_mask = 1'h1;
  assign mem_MPORT_221_en = reset;
  assign mem_MPORT_222_data = 2'h0;
  assign mem_MPORT_222_addr = 9'hde;
  assign mem_MPORT_222_mask = 1'h1;
  assign mem_MPORT_222_en = reset;
  assign mem_MPORT_223_data = 2'h0;
  assign mem_MPORT_223_addr = 9'hdf;
  assign mem_MPORT_223_mask = 1'h1;
  assign mem_MPORT_223_en = reset;
  assign mem_MPORT_224_data = 2'h0;
  assign mem_MPORT_224_addr = 9'he0;
  assign mem_MPORT_224_mask = 1'h1;
  assign mem_MPORT_224_en = reset;
  assign mem_MPORT_225_data = 2'h0;
  assign mem_MPORT_225_addr = 9'he1;
  assign mem_MPORT_225_mask = 1'h1;
  assign mem_MPORT_225_en = reset;
  assign mem_MPORT_226_data = 2'h0;
  assign mem_MPORT_226_addr = 9'he2;
  assign mem_MPORT_226_mask = 1'h1;
  assign mem_MPORT_226_en = reset;
  assign mem_MPORT_227_data = 2'h0;
  assign mem_MPORT_227_addr = 9'he3;
  assign mem_MPORT_227_mask = 1'h1;
  assign mem_MPORT_227_en = reset;
  assign mem_MPORT_228_data = 2'h0;
  assign mem_MPORT_228_addr = 9'he4;
  assign mem_MPORT_228_mask = 1'h1;
  assign mem_MPORT_228_en = reset;
  assign mem_MPORT_229_data = 2'h0;
  assign mem_MPORT_229_addr = 9'he5;
  assign mem_MPORT_229_mask = 1'h1;
  assign mem_MPORT_229_en = reset;
  assign mem_MPORT_230_data = 2'h0;
  assign mem_MPORT_230_addr = 9'he6;
  assign mem_MPORT_230_mask = 1'h1;
  assign mem_MPORT_230_en = reset;
  assign mem_MPORT_231_data = 2'h0;
  assign mem_MPORT_231_addr = 9'he7;
  assign mem_MPORT_231_mask = 1'h1;
  assign mem_MPORT_231_en = reset;
  assign mem_MPORT_232_data = 2'h0;
  assign mem_MPORT_232_addr = 9'he8;
  assign mem_MPORT_232_mask = 1'h1;
  assign mem_MPORT_232_en = reset;
  assign mem_MPORT_233_data = 2'h0;
  assign mem_MPORT_233_addr = 9'he9;
  assign mem_MPORT_233_mask = 1'h1;
  assign mem_MPORT_233_en = reset;
  assign mem_MPORT_234_data = 2'h0;
  assign mem_MPORT_234_addr = 9'hea;
  assign mem_MPORT_234_mask = 1'h1;
  assign mem_MPORT_234_en = reset;
  assign mem_MPORT_235_data = 2'h0;
  assign mem_MPORT_235_addr = 9'heb;
  assign mem_MPORT_235_mask = 1'h1;
  assign mem_MPORT_235_en = reset;
  assign mem_MPORT_236_data = 2'h0;
  assign mem_MPORT_236_addr = 9'hec;
  assign mem_MPORT_236_mask = 1'h1;
  assign mem_MPORT_236_en = reset;
  assign mem_MPORT_237_data = 2'h0;
  assign mem_MPORT_237_addr = 9'hed;
  assign mem_MPORT_237_mask = 1'h1;
  assign mem_MPORT_237_en = reset;
  assign mem_MPORT_238_data = 2'h0;
  assign mem_MPORT_238_addr = 9'hee;
  assign mem_MPORT_238_mask = 1'h1;
  assign mem_MPORT_238_en = reset;
  assign mem_MPORT_239_data = 2'h0;
  assign mem_MPORT_239_addr = 9'hef;
  assign mem_MPORT_239_mask = 1'h1;
  assign mem_MPORT_239_en = reset;
  assign mem_MPORT_240_data = 2'h0;
  assign mem_MPORT_240_addr = 9'hf0;
  assign mem_MPORT_240_mask = 1'h1;
  assign mem_MPORT_240_en = reset;
  assign mem_MPORT_241_data = 2'h0;
  assign mem_MPORT_241_addr = 9'hf1;
  assign mem_MPORT_241_mask = 1'h1;
  assign mem_MPORT_241_en = reset;
  assign mem_MPORT_242_data = 2'h0;
  assign mem_MPORT_242_addr = 9'hf2;
  assign mem_MPORT_242_mask = 1'h1;
  assign mem_MPORT_242_en = reset;
  assign mem_MPORT_243_data = 2'h0;
  assign mem_MPORT_243_addr = 9'hf3;
  assign mem_MPORT_243_mask = 1'h1;
  assign mem_MPORT_243_en = reset;
  assign mem_MPORT_244_data = 2'h0;
  assign mem_MPORT_244_addr = 9'hf4;
  assign mem_MPORT_244_mask = 1'h1;
  assign mem_MPORT_244_en = reset;
  assign mem_MPORT_245_data = 2'h0;
  assign mem_MPORT_245_addr = 9'hf5;
  assign mem_MPORT_245_mask = 1'h1;
  assign mem_MPORT_245_en = reset;
  assign mem_MPORT_246_data = 2'h0;
  assign mem_MPORT_246_addr = 9'hf6;
  assign mem_MPORT_246_mask = 1'h1;
  assign mem_MPORT_246_en = reset;
  assign mem_MPORT_247_data = 2'h0;
  assign mem_MPORT_247_addr = 9'hf7;
  assign mem_MPORT_247_mask = 1'h1;
  assign mem_MPORT_247_en = reset;
  assign mem_MPORT_248_data = 2'h0;
  assign mem_MPORT_248_addr = 9'hf8;
  assign mem_MPORT_248_mask = 1'h1;
  assign mem_MPORT_248_en = reset;
  assign mem_MPORT_249_data = 2'h0;
  assign mem_MPORT_249_addr = 9'hf9;
  assign mem_MPORT_249_mask = 1'h1;
  assign mem_MPORT_249_en = reset;
  assign mem_MPORT_250_data = 2'h0;
  assign mem_MPORT_250_addr = 9'hfa;
  assign mem_MPORT_250_mask = 1'h1;
  assign mem_MPORT_250_en = reset;
  assign mem_MPORT_251_data = 2'h0;
  assign mem_MPORT_251_addr = 9'hfb;
  assign mem_MPORT_251_mask = 1'h1;
  assign mem_MPORT_251_en = reset;
  assign mem_MPORT_252_data = 2'h0;
  assign mem_MPORT_252_addr = 9'hfc;
  assign mem_MPORT_252_mask = 1'h1;
  assign mem_MPORT_252_en = reset;
  assign mem_MPORT_253_data = 2'h0;
  assign mem_MPORT_253_addr = 9'hfd;
  assign mem_MPORT_253_mask = 1'h1;
  assign mem_MPORT_253_en = reset;
  assign mem_MPORT_254_data = 2'h0;
  assign mem_MPORT_254_addr = 9'hfe;
  assign mem_MPORT_254_mask = 1'h1;
  assign mem_MPORT_254_en = reset;
  assign mem_MPORT_255_data = 2'h0;
  assign mem_MPORT_255_addr = 9'hff;
  assign mem_MPORT_255_mask = 1'h1;
  assign mem_MPORT_255_en = reset;
  assign mem_MPORT_256_data = 2'h0;
  assign mem_MPORT_256_addr = 9'h100;
  assign mem_MPORT_256_mask = 1'h1;
  assign mem_MPORT_256_en = reset;
  assign mem_MPORT_257_data = 2'h0;
  assign mem_MPORT_257_addr = 9'h101;
  assign mem_MPORT_257_mask = 1'h1;
  assign mem_MPORT_257_en = reset;
  assign mem_MPORT_258_data = 2'h0;
  assign mem_MPORT_258_addr = 9'h102;
  assign mem_MPORT_258_mask = 1'h1;
  assign mem_MPORT_258_en = reset;
  assign mem_MPORT_259_data = 2'h0;
  assign mem_MPORT_259_addr = 9'h103;
  assign mem_MPORT_259_mask = 1'h1;
  assign mem_MPORT_259_en = reset;
  assign mem_MPORT_260_data = 2'h0;
  assign mem_MPORT_260_addr = 9'h104;
  assign mem_MPORT_260_mask = 1'h1;
  assign mem_MPORT_260_en = reset;
  assign mem_MPORT_261_data = 2'h0;
  assign mem_MPORT_261_addr = 9'h105;
  assign mem_MPORT_261_mask = 1'h1;
  assign mem_MPORT_261_en = reset;
  assign mem_MPORT_262_data = 2'h0;
  assign mem_MPORT_262_addr = 9'h106;
  assign mem_MPORT_262_mask = 1'h1;
  assign mem_MPORT_262_en = reset;
  assign mem_MPORT_263_data = 2'h0;
  assign mem_MPORT_263_addr = 9'h107;
  assign mem_MPORT_263_mask = 1'h1;
  assign mem_MPORT_263_en = reset;
  assign mem_MPORT_264_data = 2'h0;
  assign mem_MPORT_264_addr = 9'h108;
  assign mem_MPORT_264_mask = 1'h1;
  assign mem_MPORT_264_en = reset;
  assign mem_MPORT_265_data = 2'h0;
  assign mem_MPORT_265_addr = 9'h109;
  assign mem_MPORT_265_mask = 1'h1;
  assign mem_MPORT_265_en = reset;
  assign mem_MPORT_266_data = 2'h0;
  assign mem_MPORT_266_addr = 9'h10a;
  assign mem_MPORT_266_mask = 1'h1;
  assign mem_MPORT_266_en = reset;
  assign mem_MPORT_267_data = 2'h0;
  assign mem_MPORT_267_addr = 9'h10b;
  assign mem_MPORT_267_mask = 1'h1;
  assign mem_MPORT_267_en = reset;
  assign mem_MPORT_268_data = 2'h0;
  assign mem_MPORT_268_addr = 9'h10c;
  assign mem_MPORT_268_mask = 1'h1;
  assign mem_MPORT_268_en = reset;
  assign mem_MPORT_269_data = 2'h0;
  assign mem_MPORT_269_addr = 9'h10d;
  assign mem_MPORT_269_mask = 1'h1;
  assign mem_MPORT_269_en = reset;
  assign mem_MPORT_270_data = 2'h0;
  assign mem_MPORT_270_addr = 9'h10e;
  assign mem_MPORT_270_mask = 1'h1;
  assign mem_MPORT_270_en = reset;
  assign mem_MPORT_271_data = 2'h0;
  assign mem_MPORT_271_addr = 9'h10f;
  assign mem_MPORT_271_mask = 1'h1;
  assign mem_MPORT_271_en = reset;
  assign mem_MPORT_272_data = 2'h0;
  assign mem_MPORT_272_addr = 9'h110;
  assign mem_MPORT_272_mask = 1'h1;
  assign mem_MPORT_272_en = reset;
  assign mem_MPORT_273_data = 2'h0;
  assign mem_MPORT_273_addr = 9'h111;
  assign mem_MPORT_273_mask = 1'h1;
  assign mem_MPORT_273_en = reset;
  assign mem_MPORT_274_data = 2'h0;
  assign mem_MPORT_274_addr = 9'h112;
  assign mem_MPORT_274_mask = 1'h1;
  assign mem_MPORT_274_en = reset;
  assign mem_MPORT_275_data = 2'h0;
  assign mem_MPORT_275_addr = 9'h113;
  assign mem_MPORT_275_mask = 1'h1;
  assign mem_MPORT_275_en = reset;
  assign mem_MPORT_276_data = 2'h0;
  assign mem_MPORT_276_addr = 9'h114;
  assign mem_MPORT_276_mask = 1'h1;
  assign mem_MPORT_276_en = reset;
  assign mem_MPORT_277_data = 2'h0;
  assign mem_MPORT_277_addr = 9'h115;
  assign mem_MPORT_277_mask = 1'h1;
  assign mem_MPORT_277_en = reset;
  assign mem_MPORT_278_data = 2'h0;
  assign mem_MPORT_278_addr = 9'h116;
  assign mem_MPORT_278_mask = 1'h1;
  assign mem_MPORT_278_en = reset;
  assign mem_MPORT_279_data = 2'h0;
  assign mem_MPORT_279_addr = 9'h117;
  assign mem_MPORT_279_mask = 1'h1;
  assign mem_MPORT_279_en = reset;
  assign mem_MPORT_280_data = 2'h0;
  assign mem_MPORT_280_addr = 9'h118;
  assign mem_MPORT_280_mask = 1'h1;
  assign mem_MPORT_280_en = reset;
  assign mem_MPORT_281_data = 2'h0;
  assign mem_MPORT_281_addr = 9'h119;
  assign mem_MPORT_281_mask = 1'h1;
  assign mem_MPORT_281_en = reset;
  assign mem_MPORT_282_data = 2'h0;
  assign mem_MPORT_282_addr = 9'h11a;
  assign mem_MPORT_282_mask = 1'h1;
  assign mem_MPORT_282_en = reset;
  assign mem_MPORT_283_data = 2'h0;
  assign mem_MPORT_283_addr = 9'h11b;
  assign mem_MPORT_283_mask = 1'h1;
  assign mem_MPORT_283_en = reset;
  assign mem_MPORT_284_data = 2'h0;
  assign mem_MPORT_284_addr = 9'h11c;
  assign mem_MPORT_284_mask = 1'h1;
  assign mem_MPORT_284_en = reset;
  assign mem_MPORT_285_data = 2'h0;
  assign mem_MPORT_285_addr = 9'h11d;
  assign mem_MPORT_285_mask = 1'h1;
  assign mem_MPORT_285_en = reset;
  assign mem_MPORT_286_data = 2'h0;
  assign mem_MPORT_286_addr = 9'h11e;
  assign mem_MPORT_286_mask = 1'h1;
  assign mem_MPORT_286_en = reset;
  assign mem_MPORT_287_data = 2'h0;
  assign mem_MPORT_287_addr = 9'h11f;
  assign mem_MPORT_287_mask = 1'h1;
  assign mem_MPORT_287_en = reset;
  assign mem_MPORT_288_data = 2'h0;
  assign mem_MPORT_288_addr = 9'h120;
  assign mem_MPORT_288_mask = 1'h1;
  assign mem_MPORT_288_en = reset;
  assign mem_MPORT_289_data = 2'h0;
  assign mem_MPORT_289_addr = 9'h121;
  assign mem_MPORT_289_mask = 1'h1;
  assign mem_MPORT_289_en = reset;
  assign mem_MPORT_290_data = 2'h0;
  assign mem_MPORT_290_addr = 9'h122;
  assign mem_MPORT_290_mask = 1'h1;
  assign mem_MPORT_290_en = reset;
  assign mem_MPORT_291_data = 2'h0;
  assign mem_MPORT_291_addr = 9'h123;
  assign mem_MPORT_291_mask = 1'h1;
  assign mem_MPORT_291_en = reset;
  assign mem_MPORT_292_data = 2'h0;
  assign mem_MPORT_292_addr = 9'h124;
  assign mem_MPORT_292_mask = 1'h1;
  assign mem_MPORT_292_en = reset;
  assign mem_MPORT_293_data = 2'h0;
  assign mem_MPORT_293_addr = 9'h125;
  assign mem_MPORT_293_mask = 1'h1;
  assign mem_MPORT_293_en = reset;
  assign mem_MPORT_294_data = 2'h0;
  assign mem_MPORT_294_addr = 9'h126;
  assign mem_MPORT_294_mask = 1'h1;
  assign mem_MPORT_294_en = reset;
  assign mem_MPORT_295_data = 2'h0;
  assign mem_MPORT_295_addr = 9'h127;
  assign mem_MPORT_295_mask = 1'h1;
  assign mem_MPORT_295_en = reset;
  assign mem_MPORT_296_data = 2'h0;
  assign mem_MPORT_296_addr = 9'h128;
  assign mem_MPORT_296_mask = 1'h1;
  assign mem_MPORT_296_en = reset;
  assign mem_MPORT_297_data = 2'h0;
  assign mem_MPORT_297_addr = 9'h129;
  assign mem_MPORT_297_mask = 1'h1;
  assign mem_MPORT_297_en = reset;
  assign mem_MPORT_298_data = 2'h0;
  assign mem_MPORT_298_addr = 9'h12a;
  assign mem_MPORT_298_mask = 1'h1;
  assign mem_MPORT_298_en = reset;
  assign mem_MPORT_299_data = 2'h0;
  assign mem_MPORT_299_addr = 9'h12b;
  assign mem_MPORT_299_mask = 1'h1;
  assign mem_MPORT_299_en = reset;
  assign mem_MPORT_300_data = 2'h0;
  assign mem_MPORT_300_addr = 9'h12c;
  assign mem_MPORT_300_mask = 1'h1;
  assign mem_MPORT_300_en = reset;
  assign mem_MPORT_301_data = 2'h0;
  assign mem_MPORT_301_addr = 9'h12d;
  assign mem_MPORT_301_mask = 1'h1;
  assign mem_MPORT_301_en = reset;
  assign mem_MPORT_302_data = 2'h0;
  assign mem_MPORT_302_addr = 9'h12e;
  assign mem_MPORT_302_mask = 1'h1;
  assign mem_MPORT_302_en = reset;
  assign mem_MPORT_303_data = 2'h0;
  assign mem_MPORT_303_addr = 9'h12f;
  assign mem_MPORT_303_mask = 1'h1;
  assign mem_MPORT_303_en = reset;
  assign mem_MPORT_304_data = 2'h0;
  assign mem_MPORT_304_addr = 9'h130;
  assign mem_MPORT_304_mask = 1'h1;
  assign mem_MPORT_304_en = reset;
  assign mem_MPORT_305_data = 2'h0;
  assign mem_MPORT_305_addr = 9'h131;
  assign mem_MPORT_305_mask = 1'h1;
  assign mem_MPORT_305_en = reset;
  assign mem_MPORT_306_data = 2'h0;
  assign mem_MPORT_306_addr = 9'h132;
  assign mem_MPORT_306_mask = 1'h1;
  assign mem_MPORT_306_en = reset;
  assign mem_MPORT_307_data = 2'h0;
  assign mem_MPORT_307_addr = 9'h133;
  assign mem_MPORT_307_mask = 1'h1;
  assign mem_MPORT_307_en = reset;
  assign mem_MPORT_308_data = 2'h0;
  assign mem_MPORT_308_addr = 9'h134;
  assign mem_MPORT_308_mask = 1'h1;
  assign mem_MPORT_308_en = reset;
  assign mem_MPORT_309_data = 2'h0;
  assign mem_MPORT_309_addr = 9'h135;
  assign mem_MPORT_309_mask = 1'h1;
  assign mem_MPORT_309_en = reset;
  assign mem_MPORT_310_data = 2'h0;
  assign mem_MPORT_310_addr = 9'h136;
  assign mem_MPORT_310_mask = 1'h1;
  assign mem_MPORT_310_en = reset;
  assign mem_MPORT_311_data = 2'h0;
  assign mem_MPORT_311_addr = 9'h137;
  assign mem_MPORT_311_mask = 1'h1;
  assign mem_MPORT_311_en = reset;
  assign mem_MPORT_312_data = 2'h0;
  assign mem_MPORT_312_addr = 9'h138;
  assign mem_MPORT_312_mask = 1'h1;
  assign mem_MPORT_312_en = reset;
  assign mem_MPORT_313_data = 2'h0;
  assign mem_MPORT_313_addr = 9'h139;
  assign mem_MPORT_313_mask = 1'h1;
  assign mem_MPORT_313_en = reset;
  assign mem_MPORT_314_data = 2'h0;
  assign mem_MPORT_314_addr = 9'h13a;
  assign mem_MPORT_314_mask = 1'h1;
  assign mem_MPORT_314_en = reset;
  assign mem_MPORT_315_data = 2'h0;
  assign mem_MPORT_315_addr = 9'h13b;
  assign mem_MPORT_315_mask = 1'h1;
  assign mem_MPORT_315_en = reset;
  assign mem_MPORT_316_data = 2'h0;
  assign mem_MPORT_316_addr = 9'h13c;
  assign mem_MPORT_316_mask = 1'h1;
  assign mem_MPORT_316_en = reset;
  assign mem_MPORT_317_data = 2'h0;
  assign mem_MPORT_317_addr = 9'h13d;
  assign mem_MPORT_317_mask = 1'h1;
  assign mem_MPORT_317_en = reset;
  assign mem_MPORT_318_data = 2'h0;
  assign mem_MPORT_318_addr = 9'h13e;
  assign mem_MPORT_318_mask = 1'h1;
  assign mem_MPORT_318_en = reset;
  assign mem_MPORT_319_data = 2'h0;
  assign mem_MPORT_319_addr = 9'h13f;
  assign mem_MPORT_319_mask = 1'h1;
  assign mem_MPORT_319_en = reset;
  assign mem_MPORT_320_data = 2'h0;
  assign mem_MPORT_320_addr = 9'h140;
  assign mem_MPORT_320_mask = 1'h1;
  assign mem_MPORT_320_en = reset;
  assign mem_MPORT_321_data = 2'h0;
  assign mem_MPORT_321_addr = 9'h141;
  assign mem_MPORT_321_mask = 1'h1;
  assign mem_MPORT_321_en = reset;
  assign mem_MPORT_322_data = 2'h0;
  assign mem_MPORT_322_addr = 9'h142;
  assign mem_MPORT_322_mask = 1'h1;
  assign mem_MPORT_322_en = reset;
  assign mem_MPORT_323_data = 2'h0;
  assign mem_MPORT_323_addr = 9'h143;
  assign mem_MPORT_323_mask = 1'h1;
  assign mem_MPORT_323_en = reset;
  assign mem_MPORT_324_data = 2'h0;
  assign mem_MPORT_324_addr = 9'h144;
  assign mem_MPORT_324_mask = 1'h1;
  assign mem_MPORT_324_en = reset;
  assign mem_MPORT_325_data = 2'h0;
  assign mem_MPORT_325_addr = 9'h145;
  assign mem_MPORT_325_mask = 1'h1;
  assign mem_MPORT_325_en = reset;
  assign mem_MPORT_326_data = 2'h0;
  assign mem_MPORT_326_addr = 9'h146;
  assign mem_MPORT_326_mask = 1'h1;
  assign mem_MPORT_326_en = reset;
  assign mem_MPORT_327_data = 2'h0;
  assign mem_MPORT_327_addr = 9'h147;
  assign mem_MPORT_327_mask = 1'h1;
  assign mem_MPORT_327_en = reset;
  assign mem_MPORT_328_data = 2'h0;
  assign mem_MPORT_328_addr = 9'h148;
  assign mem_MPORT_328_mask = 1'h1;
  assign mem_MPORT_328_en = reset;
  assign mem_MPORT_329_data = 2'h0;
  assign mem_MPORT_329_addr = 9'h149;
  assign mem_MPORT_329_mask = 1'h1;
  assign mem_MPORT_329_en = reset;
  assign mem_MPORT_330_data = 2'h0;
  assign mem_MPORT_330_addr = 9'h14a;
  assign mem_MPORT_330_mask = 1'h1;
  assign mem_MPORT_330_en = reset;
  assign mem_MPORT_331_data = 2'h0;
  assign mem_MPORT_331_addr = 9'h14b;
  assign mem_MPORT_331_mask = 1'h1;
  assign mem_MPORT_331_en = reset;
  assign mem_MPORT_332_data = 2'h0;
  assign mem_MPORT_332_addr = 9'h14c;
  assign mem_MPORT_332_mask = 1'h1;
  assign mem_MPORT_332_en = reset;
  assign mem_MPORT_333_data = 2'h0;
  assign mem_MPORT_333_addr = 9'h14d;
  assign mem_MPORT_333_mask = 1'h1;
  assign mem_MPORT_333_en = reset;
  assign mem_MPORT_334_data = 2'h0;
  assign mem_MPORT_334_addr = 9'h14e;
  assign mem_MPORT_334_mask = 1'h1;
  assign mem_MPORT_334_en = reset;
  assign mem_MPORT_335_data = 2'h0;
  assign mem_MPORT_335_addr = 9'h14f;
  assign mem_MPORT_335_mask = 1'h1;
  assign mem_MPORT_335_en = reset;
  assign mem_MPORT_336_data = 2'h0;
  assign mem_MPORT_336_addr = 9'h150;
  assign mem_MPORT_336_mask = 1'h1;
  assign mem_MPORT_336_en = reset;
  assign mem_MPORT_337_data = 2'h0;
  assign mem_MPORT_337_addr = 9'h151;
  assign mem_MPORT_337_mask = 1'h1;
  assign mem_MPORT_337_en = reset;
  assign mem_MPORT_338_data = 2'h0;
  assign mem_MPORT_338_addr = 9'h152;
  assign mem_MPORT_338_mask = 1'h1;
  assign mem_MPORT_338_en = reset;
  assign mem_MPORT_339_data = 2'h0;
  assign mem_MPORT_339_addr = 9'h153;
  assign mem_MPORT_339_mask = 1'h1;
  assign mem_MPORT_339_en = reset;
  assign mem_MPORT_340_data = 2'h0;
  assign mem_MPORT_340_addr = 9'h154;
  assign mem_MPORT_340_mask = 1'h1;
  assign mem_MPORT_340_en = reset;
  assign mem_MPORT_341_data = 2'h0;
  assign mem_MPORT_341_addr = 9'h155;
  assign mem_MPORT_341_mask = 1'h1;
  assign mem_MPORT_341_en = reset;
  assign mem_MPORT_342_data = 2'h0;
  assign mem_MPORT_342_addr = 9'h156;
  assign mem_MPORT_342_mask = 1'h1;
  assign mem_MPORT_342_en = reset;
  assign mem_MPORT_343_data = 2'h0;
  assign mem_MPORT_343_addr = 9'h157;
  assign mem_MPORT_343_mask = 1'h1;
  assign mem_MPORT_343_en = reset;
  assign mem_MPORT_344_data = 2'h0;
  assign mem_MPORT_344_addr = 9'h158;
  assign mem_MPORT_344_mask = 1'h1;
  assign mem_MPORT_344_en = reset;
  assign mem_MPORT_345_data = 2'h0;
  assign mem_MPORT_345_addr = 9'h159;
  assign mem_MPORT_345_mask = 1'h1;
  assign mem_MPORT_345_en = reset;
  assign mem_MPORT_346_data = 2'h0;
  assign mem_MPORT_346_addr = 9'h15a;
  assign mem_MPORT_346_mask = 1'h1;
  assign mem_MPORT_346_en = reset;
  assign mem_MPORT_347_data = 2'h0;
  assign mem_MPORT_347_addr = 9'h15b;
  assign mem_MPORT_347_mask = 1'h1;
  assign mem_MPORT_347_en = reset;
  assign mem_MPORT_348_data = 2'h0;
  assign mem_MPORT_348_addr = 9'h15c;
  assign mem_MPORT_348_mask = 1'h1;
  assign mem_MPORT_348_en = reset;
  assign mem_MPORT_349_data = 2'h0;
  assign mem_MPORT_349_addr = 9'h15d;
  assign mem_MPORT_349_mask = 1'h1;
  assign mem_MPORT_349_en = reset;
  assign mem_MPORT_350_data = 2'h0;
  assign mem_MPORT_350_addr = 9'h15e;
  assign mem_MPORT_350_mask = 1'h1;
  assign mem_MPORT_350_en = reset;
  assign mem_MPORT_351_data = 2'h0;
  assign mem_MPORT_351_addr = 9'h15f;
  assign mem_MPORT_351_mask = 1'h1;
  assign mem_MPORT_351_en = reset;
  assign mem_MPORT_352_data = 2'h0;
  assign mem_MPORT_352_addr = 9'h160;
  assign mem_MPORT_352_mask = 1'h1;
  assign mem_MPORT_352_en = reset;
  assign mem_MPORT_353_data = 2'h0;
  assign mem_MPORT_353_addr = 9'h161;
  assign mem_MPORT_353_mask = 1'h1;
  assign mem_MPORT_353_en = reset;
  assign mem_MPORT_354_data = 2'h0;
  assign mem_MPORT_354_addr = 9'h162;
  assign mem_MPORT_354_mask = 1'h1;
  assign mem_MPORT_354_en = reset;
  assign mem_MPORT_355_data = 2'h0;
  assign mem_MPORT_355_addr = 9'h163;
  assign mem_MPORT_355_mask = 1'h1;
  assign mem_MPORT_355_en = reset;
  assign mem_MPORT_356_data = 2'h0;
  assign mem_MPORT_356_addr = 9'h164;
  assign mem_MPORT_356_mask = 1'h1;
  assign mem_MPORT_356_en = reset;
  assign mem_MPORT_357_data = 2'h0;
  assign mem_MPORT_357_addr = 9'h165;
  assign mem_MPORT_357_mask = 1'h1;
  assign mem_MPORT_357_en = reset;
  assign mem_MPORT_358_data = 2'h0;
  assign mem_MPORT_358_addr = 9'h166;
  assign mem_MPORT_358_mask = 1'h1;
  assign mem_MPORT_358_en = reset;
  assign mem_MPORT_359_data = 2'h0;
  assign mem_MPORT_359_addr = 9'h167;
  assign mem_MPORT_359_mask = 1'h1;
  assign mem_MPORT_359_en = reset;
  assign mem_MPORT_360_data = 2'h0;
  assign mem_MPORT_360_addr = 9'h168;
  assign mem_MPORT_360_mask = 1'h1;
  assign mem_MPORT_360_en = reset;
  assign mem_MPORT_361_data = 2'h0;
  assign mem_MPORT_361_addr = 9'h169;
  assign mem_MPORT_361_mask = 1'h1;
  assign mem_MPORT_361_en = reset;
  assign mem_MPORT_362_data = 2'h0;
  assign mem_MPORT_362_addr = 9'h16a;
  assign mem_MPORT_362_mask = 1'h1;
  assign mem_MPORT_362_en = reset;
  assign mem_MPORT_363_data = 2'h0;
  assign mem_MPORT_363_addr = 9'h16b;
  assign mem_MPORT_363_mask = 1'h1;
  assign mem_MPORT_363_en = reset;
  assign mem_MPORT_364_data = 2'h0;
  assign mem_MPORT_364_addr = 9'h16c;
  assign mem_MPORT_364_mask = 1'h1;
  assign mem_MPORT_364_en = reset;
  assign mem_MPORT_365_data = 2'h0;
  assign mem_MPORT_365_addr = 9'h16d;
  assign mem_MPORT_365_mask = 1'h1;
  assign mem_MPORT_365_en = reset;
  assign mem_MPORT_366_data = 2'h0;
  assign mem_MPORT_366_addr = 9'h16e;
  assign mem_MPORT_366_mask = 1'h1;
  assign mem_MPORT_366_en = reset;
  assign mem_MPORT_367_data = 2'h0;
  assign mem_MPORT_367_addr = 9'h16f;
  assign mem_MPORT_367_mask = 1'h1;
  assign mem_MPORT_367_en = reset;
  assign mem_MPORT_368_data = 2'h0;
  assign mem_MPORT_368_addr = 9'h170;
  assign mem_MPORT_368_mask = 1'h1;
  assign mem_MPORT_368_en = reset;
  assign mem_MPORT_369_data = 2'h0;
  assign mem_MPORT_369_addr = 9'h171;
  assign mem_MPORT_369_mask = 1'h1;
  assign mem_MPORT_369_en = reset;
  assign mem_MPORT_370_data = 2'h0;
  assign mem_MPORT_370_addr = 9'h172;
  assign mem_MPORT_370_mask = 1'h1;
  assign mem_MPORT_370_en = reset;
  assign mem_MPORT_371_data = 2'h0;
  assign mem_MPORT_371_addr = 9'h173;
  assign mem_MPORT_371_mask = 1'h1;
  assign mem_MPORT_371_en = reset;
  assign mem_MPORT_372_data = 2'h0;
  assign mem_MPORT_372_addr = 9'h174;
  assign mem_MPORT_372_mask = 1'h1;
  assign mem_MPORT_372_en = reset;
  assign mem_MPORT_373_data = 2'h0;
  assign mem_MPORT_373_addr = 9'h175;
  assign mem_MPORT_373_mask = 1'h1;
  assign mem_MPORT_373_en = reset;
  assign mem_MPORT_374_data = 2'h0;
  assign mem_MPORT_374_addr = 9'h176;
  assign mem_MPORT_374_mask = 1'h1;
  assign mem_MPORT_374_en = reset;
  assign mem_MPORT_375_data = 2'h0;
  assign mem_MPORT_375_addr = 9'h177;
  assign mem_MPORT_375_mask = 1'h1;
  assign mem_MPORT_375_en = reset;
  assign mem_MPORT_376_data = 2'h0;
  assign mem_MPORT_376_addr = 9'h178;
  assign mem_MPORT_376_mask = 1'h1;
  assign mem_MPORT_376_en = reset;
  assign mem_MPORT_377_data = 2'h0;
  assign mem_MPORT_377_addr = 9'h179;
  assign mem_MPORT_377_mask = 1'h1;
  assign mem_MPORT_377_en = reset;
  assign mem_MPORT_378_data = 2'h0;
  assign mem_MPORT_378_addr = 9'h17a;
  assign mem_MPORT_378_mask = 1'h1;
  assign mem_MPORT_378_en = reset;
  assign mem_MPORT_379_data = 2'h0;
  assign mem_MPORT_379_addr = 9'h17b;
  assign mem_MPORT_379_mask = 1'h1;
  assign mem_MPORT_379_en = reset;
  assign mem_MPORT_380_data = 2'h0;
  assign mem_MPORT_380_addr = 9'h17c;
  assign mem_MPORT_380_mask = 1'h1;
  assign mem_MPORT_380_en = reset;
  assign mem_MPORT_381_data = 2'h0;
  assign mem_MPORT_381_addr = 9'h17d;
  assign mem_MPORT_381_mask = 1'h1;
  assign mem_MPORT_381_en = reset;
  assign mem_MPORT_382_data = 2'h0;
  assign mem_MPORT_382_addr = 9'h17e;
  assign mem_MPORT_382_mask = 1'h1;
  assign mem_MPORT_382_en = reset;
  assign mem_MPORT_383_data = 2'h0;
  assign mem_MPORT_383_addr = 9'h17f;
  assign mem_MPORT_383_mask = 1'h1;
  assign mem_MPORT_383_en = reset;
  assign mem_MPORT_384_data = 2'h0;
  assign mem_MPORT_384_addr = 9'h180;
  assign mem_MPORT_384_mask = 1'h1;
  assign mem_MPORT_384_en = reset;
  assign mem_MPORT_385_data = 2'h0;
  assign mem_MPORT_385_addr = 9'h181;
  assign mem_MPORT_385_mask = 1'h1;
  assign mem_MPORT_385_en = reset;
  assign mem_MPORT_386_data = 2'h0;
  assign mem_MPORT_386_addr = 9'h182;
  assign mem_MPORT_386_mask = 1'h1;
  assign mem_MPORT_386_en = reset;
  assign mem_MPORT_387_data = 2'h0;
  assign mem_MPORT_387_addr = 9'h183;
  assign mem_MPORT_387_mask = 1'h1;
  assign mem_MPORT_387_en = reset;
  assign mem_MPORT_388_data = 2'h0;
  assign mem_MPORT_388_addr = 9'h184;
  assign mem_MPORT_388_mask = 1'h1;
  assign mem_MPORT_388_en = reset;
  assign mem_MPORT_389_data = 2'h0;
  assign mem_MPORT_389_addr = 9'h185;
  assign mem_MPORT_389_mask = 1'h1;
  assign mem_MPORT_389_en = reset;
  assign mem_MPORT_390_data = 2'h0;
  assign mem_MPORT_390_addr = 9'h186;
  assign mem_MPORT_390_mask = 1'h1;
  assign mem_MPORT_390_en = reset;
  assign mem_MPORT_391_data = 2'h0;
  assign mem_MPORT_391_addr = 9'h187;
  assign mem_MPORT_391_mask = 1'h1;
  assign mem_MPORT_391_en = reset;
  assign mem_MPORT_392_data = 2'h0;
  assign mem_MPORT_392_addr = 9'h188;
  assign mem_MPORT_392_mask = 1'h1;
  assign mem_MPORT_392_en = reset;
  assign mem_MPORT_393_data = 2'h0;
  assign mem_MPORT_393_addr = 9'h189;
  assign mem_MPORT_393_mask = 1'h1;
  assign mem_MPORT_393_en = reset;
  assign mem_MPORT_394_data = 2'h0;
  assign mem_MPORT_394_addr = 9'h18a;
  assign mem_MPORT_394_mask = 1'h1;
  assign mem_MPORT_394_en = reset;
  assign mem_MPORT_395_data = 2'h0;
  assign mem_MPORT_395_addr = 9'h18b;
  assign mem_MPORT_395_mask = 1'h1;
  assign mem_MPORT_395_en = reset;
  assign mem_MPORT_396_data = 2'h0;
  assign mem_MPORT_396_addr = 9'h18c;
  assign mem_MPORT_396_mask = 1'h1;
  assign mem_MPORT_396_en = reset;
  assign mem_MPORT_397_data = 2'h0;
  assign mem_MPORT_397_addr = 9'h18d;
  assign mem_MPORT_397_mask = 1'h1;
  assign mem_MPORT_397_en = reset;
  assign mem_MPORT_398_data = 2'h0;
  assign mem_MPORT_398_addr = 9'h18e;
  assign mem_MPORT_398_mask = 1'h1;
  assign mem_MPORT_398_en = reset;
  assign mem_MPORT_399_data = 2'h0;
  assign mem_MPORT_399_addr = 9'h18f;
  assign mem_MPORT_399_mask = 1'h1;
  assign mem_MPORT_399_en = reset;
  assign mem_MPORT_400_data = 2'h0;
  assign mem_MPORT_400_addr = 9'h190;
  assign mem_MPORT_400_mask = 1'h1;
  assign mem_MPORT_400_en = reset;
  assign mem_MPORT_401_data = 2'h0;
  assign mem_MPORT_401_addr = 9'h191;
  assign mem_MPORT_401_mask = 1'h1;
  assign mem_MPORT_401_en = reset;
  assign mem_MPORT_402_data = 2'h0;
  assign mem_MPORT_402_addr = 9'h192;
  assign mem_MPORT_402_mask = 1'h1;
  assign mem_MPORT_402_en = reset;
  assign mem_MPORT_403_data = 2'h0;
  assign mem_MPORT_403_addr = 9'h193;
  assign mem_MPORT_403_mask = 1'h1;
  assign mem_MPORT_403_en = reset;
  assign mem_MPORT_404_data = 2'h0;
  assign mem_MPORT_404_addr = 9'h194;
  assign mem_MPORT_404_mask = 1'h1;
  assign mem_MPORT_404_en = reset;
  assign mem_MPORT_405_data = 2'h0;
  assign mem_MPORT_405_addr = 9'h195;
  assign mem_MPORT_405_mask = 1'h1;
  assign mem_MPORT_405_en = reset;
  assign mem_MPORT_406_data = 2'h0;
  assign mem_MPORT_406_addr = 9'h196;
  assign mem_MPORT_406_mask = 1'h1;
  assign mem_MPORT_406_en = reset;
  assign mem_MPORT_407_data = 2'h0;
  assign mem_MPORT_407_addr = 9'h197;
  assign mem_MPORT_407_mask = 1'h1;
  assign mem_MPORT_407_en = reset;
  assign mem_MPORT_408_data = 2'h0;
  assign mem_MPORT_408_addr = 9'h198;
  assign mem_MPORT_408_mask = 1'h1;
  assign mem_MPORT_408_en = reset;
  assign mem_MPORT_409_data = 2'h0;
  assign mem_MPORT_409_addr = 9'h199;
  assign mem_MPORT_409_mask = 1'h1;
  assign mem_MPORT_409_en = reset;
  assign mem_MPORT_410_data = 2'h0;
  assign mem_MPORT_410_addr = 9'h19a;
  assign mem_MPORT_410_mask = 1'h1;
  assign mem_MPORT_410_en = reset;
  assign mem_MPORT_411_data = 2'h0;
  assign mem_MPORT_411_addr = 9'h19b;
  assign mem_MPORT_411_mask = 1'h1;
  assign mem_MPORT_411_en = reset;
  assign mem_MPORT_412_data = 2'h0;
  assign mem_MPORT_412_addr = 9'h19c;
  assign mem_MPORT_412_mask = 1'h1;
  assign mem_MPORT_412_en = reset;
  assign mem_MPORT_413_data = 2'h0;
  assign mem_MPORT_413_addr = 9'h19d;
  assign mem_MPORT_413_mask = 1'h1;
  assign mem_MPORT_413_en = reset;
  assign mem_MPORT_414_data = 2'h0;
  assign mem_MPORT_414_addr = 9'h19e;
  assign mem_MPORT_414_mask = 1'h1;
  assign mem_MPORT_414_en = reset;
  assign mem_MPORT_415_data = 2'h0;
  assign mem_MPORT_415_addr = 9'h19f;
  assign mem_MPORT_415_mask = 1'h1;
  assign mem_MPORT_415_en = reset;
  assign mem_MPORT_416_data = 2'h0;
  assign mem_MPORT_416_addr = 9'h1a0;
  assign mem_MPORT_416_mask = 1'h1;
  assign mem_MPORT_416_en = reset;
  assign mem_MPORT_417_data = 2'h0;
  assign mem_MPORT_417_addr = 9'h1a1;
  assign mem_MPORT_417_mask = 1'h1;
  assign mem_MPORT_417_en = reset;
  assign mem_MPORT_418_data = 2'h0;
  assign mem_MPORT_418_addr = 9'h1a2;
  assign mem_MPORT_418_mask = 1'h1;
  assign mem_MPORT_418_en = reset;
  assign mem_MPORT_419_data = 2'h0;
  assign mem_MPORT_419_addr = 9'h1a3;
  assign mem_MPORT_419_mask = 1'h1;
  assign mem_MPORT_419_en = reset;
  assign mem_MPORT_420_data = 2'h0;
  assign mem_MPORT_420_addr = 9'h1a4;
  assign mem_MPORT_420_mask = 1'h1;
  assign mem_MPORT_420_en = reset;
  assign mem_MPORT_421_data = 2'h0;
  assign mem_MPORT_421_addr = 9'h1a5;
  assign mem_MPORT_421_mask = 1'h1;
  assign mem_MPORT_421_en = reset;
  assign mem_MPORT_422_data = 2'h0;
  assign mem_MPORT_422_addr = 9'h1a6;
  assign mem_MPORT_422_mask = 1'h1;
  assign mem_MPORT_422_en = reset;
  assign mem_MPORT_423_data = 2'h0;
  assign mem_MPORT_423_addr = 9'h1a7;
  assign mem_MPORT_423_mask = 1'h1;
  assign mem_MPORT_423_en = reset;
  assign mem_MPORT_424_data = 2'h0;
  assign mem_MPORT_424_addr = 9'h1a8;
  assign mem_MPORT_424_mask = 1'h1;
  assign mem_MPORT_424_en = reset;
  assign mem_MPORT_425_data = 2'h0;
  assign mem_MPORT_425_addr = 9'h1a9;
  assign mem_MPORT_425_mask = 1'h1;
  assign mem_MPORT_425_en = reset;
  assign mem_MPORT_426_data = 2'h0;
  assign mem_MPORT_426_addr = 9'h1aa;
  assign mem_MPORT_426_mask = 1'h1;
  assign mem_MPORT_426_en = reset;
  assign mem_MPORT_427_data = 2'h0;
  assign mem_MPORT_427_addr = 9'h1ab;
  assign mem_MPORT_427_mask = 1'h1;
  assign mem_MPORT_427_en = reset;
  assign mem_MPORT_428_data = 2'h0;
  assign mem_MPORT_428_addr = 9'h1ac;
  assign mem_MPORT_428_mask = 1'h1;
  assign mem_MPORT_428_en = reset;
  assign mem_MPORT_429_data = 2'h0;
  assign mem_MPORT_429_addr = 9'h1ad;
  assign mem_MPORT_429_mask = 1'h1;
  assign mem_MPORT_429_en = reset;
  assign mem_MPORT_430_data = 2'h0;
  assign mem_MPORT_430_addr = 9'h1ae;
  assign mem_MPORT_430_mask = 1'h1;
  assign mem_MPORT_430_en = reset;
  assign mem_MPORT_431_data = 2'h0;
  assign mem_MPORT_431_addr = 9'h1af;
  assign mem_MPORT_431_mask = 1'h1;
  assign mem_MPORT_431_en = reset;
  assign mem_MPORT_432_data = 2'h0;
  assign mem_MPORT_432_addr = 9'h1b0;
  assign mem_MPORT_432_mask = 1'h1;
  assign mem_MPORT_432_en = reset;
  assign mem_MPORT_433_data = 2'h0;
  assign mem_MPORT_433_addr = 9'h1b1;
  assign mem_MPORT_433_mask = 1'h1;
  assign mem_MPORT_433_en = reset;
  assign mem_MPORT_434_data = 2'h0;
  assign mem_MPORT_434_addr = 9'h1b2;
  assign mem_MPORT_434_mask = 1'h1;
  assign mem_MPORT_434_en = reset;
  assign mem_MPORT_435_data = 2'h0;
  assign mem_MPORT_435_addr = 9'h1b3;
  assign mem_MPORT_435_mask = 1'h1;
  assign mem_MPORT_435_en = reset;
  assign mem_MPORT_436_data = 2'h0;
  assign mem_MPORT_436_addr = 9'h1b4;
  assign mem_MPORT_436_mask = 1'h1;
  assign mem_MPORT_436_en = reset;
  assign mem_MPORT_437_data = 2'h0;
  assign mem_MPORT_437_addr = 9'h1b5;
  assign mem_MPORT_437_mask = 1'h1;
  assign mem_MPORT_437_en = reset;
  assign mem_MPORT_438_data = 2'h0;
  assign mem_MPORT_438_addr = 9'h1b6;
  assign mem_MPORT_438_mask = 1'h1;
  assign mem_MPORT_438_en = reset;
  assign mem_MPORT_439_data = 2'h0;
  assign mem_MPORT_439_addr = 9'h1b7;
  assign mem_MPORT_439_mask = 1'h1;
  assign mem_MPORT_439_en = reset;
  assign mem_MPORT_440_data = 2'h0;
  assign mem_MPORT_440_addr = 9'h1b8;
  assign mem_MPORT_440_mask = 1'h1;
  assign mem_MPORT_440_en = reset;
  assign mem_MPORT_441_data = 2'h0;
  assign mem_MPORT_441_addr = 9'h1b9;
  assign mem_MPORT_441_mask = 1'h1;
  assign mem_MPORT_441_en = reset;
  assign mem_MPORT_442_data = 2'h0;
  assign mem_MPORT_442_addr = 9'h1ba;
  assign mem_MPORT_442_mask = 1'h1;
  assign mem_MPORT_442_en = reset;
  assign mem_MPORT_443_data = 2'h0;
  assign mem_MPORT_443_addr = 9'h1bb;
  assign mem_MPORT_443_mask = 1'h1;
  assign mem_MPORT_443_en = reset;
  assign mem_MPORT_444_data = 2'h0;
  assign mem_MPORT_444_addr = 9'h1bc;
  assign mem_MPORT_444_mask = 1'h1;
  assign mem_MPORT_444_en = reset;
  assign mem_MPORT_445_data = 2'h0;
  assign mem_MPORT_445_addr = 9'h1bd;
  assign mem_MPORT_445_mask = 1'h1;
  assign mem_MPORT_445_en = reset;
  assign mem_MPORT_446_data = 2'h0;
  assign mem_MPORT_446_addr = 9'h1be;
  assign mem_MPORT_446_mask = 1'h1;
  assign mem_MPORT_446_en = reset;
  assign mem_MPORT_447_data = 2'h0;
  assign mem_MPORT_447_addr = 9'h1bf;
  assign mem_MPORT_447_mask = 1'h1;
  assign mem_MPORT_447_en = reset;
  assign mem_MPORT_448_data = 2'h0;
  assign mem_MPORT_448_addr = 9'h1c0;
  assign mem_MPORT_448_mask = 1'h1;
  assign mem_MPORT_448_en = reset;
  assign mem_MPORT_449_data = 2'h0;
  assign mem_MPORT_449_addr = 9'h1c1;
  assign mem_MPORT_449_mask = 1'h1;
  assign mem_MPORT_449_en = reset;
  assign mem_MPORT_450_data = 2'h0;
  assign mem_MPORT_450_addr = 9'h1c2;
  assign mem_MPORT_450_mask = 1'h1;
  assign mem_MPORT_450_en = reset;
  assign mem_MPORT_451_data = 2'h0;
  assign mem_MPORT_451_addr = 9'h1c3;
  assign mem_MPORT_451_mask = 1'h1;
  assign mem_MPORT_451_en = reset;
  assign mem_MPORT_452_data = 2'h0;
  assign mem_MPORT_452_addr = 9'h1c4;
  assign mem_MPORT_452_mask = 1'h1;
  assign mem_MPORT_452_en = reset;
  assign mem_MPORT_453_data = 2'h0;
  assign mem_MPORT_453_addr = 9'h1c5;
  assign mem_MPORT_453_mask = 1'h1;
  assign mem_MPORT_453_en = reset;
  assign mem_MPORT_454_data = 2'h0;
  assign mem_MPORT_454_addr = 9'h1c6;
  assign mem_MPORT_454_mask = 1'h1;
  assign mem_MPORT_454_en = reset;
  assign mem_MPORT_455_data = 2'h0;
  assign mem_MPORT_455_addr = 9'h1c7;
  assign mem_MPORT_455_mask = 1'h1;
  assign mem_MPORT_455_en = reset;
  assign mem_MPORT_456_data = 2'h0;
  assign mem_MPORT_456_addr = 9'h1c8;
  assign mem_MPORT_456_mask = 1'h1;
  assign mem_MPORT_456_en = reset;
  assign mem_MPORT_457_data = 2'h0;
  assign mem_MPORT_457_addr = 9'h1c9;
  assign mem_MPORT_457_mask = 1'h1;
  assign mem_MPORT_457_en = reset;
  assign mem_MPORT_458_data = 2'h0;
  assign mem_MPORT_458_addr = 9'h1ca;
  assign mem_MPORT_458_mask = 1'h1;
  assign mem_MPORT_458_en = reset;
  assign mem_MPORT_459_data = 2'h0;
  assign mem_MPORT_459_addr = 9'h1cb;
  assign mem_MPORT_459_mask = 1'h1;
  assign mem_MPORT_459_en = reset;
  assign mem_MPORT_460_data = 2'h0;
  assign mem_MPORT_460_addr = 9'h1cc;
  assign mem_MPORT_460_mask = 1'h1;
  assign mem_MPORT_460_en = reset;
  assign mem_MPORT_461_data = 2'h0;
  assign mem_MPORT_461_addr = 9'h1cd;
  assign mem_MPORT_461_mask = 1'h1;
  assign mem_MPORT_461_en = reset;
  assign mem_MPORT_462_data = 2'h0;
  assign mem_MPORT_462_addr = 9'h1ce;
  assign mem_MPORT_462_mask = 1'h1;
  assign mem_MPORT_462_en = reset;
  assign mem_MPORT_463_data = 2'h0;
  assign mem_MPORT_463_addr = 9'h1cf;
  assign mem_MPORT_463_mask = 1'h1;
  assign mem_MPORT_463_en = reset;
  assign mem_MPORT_464_data = 2'h0;
  assign mem_MPORT_464_addr = 9'h1d0;
  assign mem_MPORT_464_mask = 1'h1;
  assign mem_MPORT_464_en = reset;
  assign mem_MPORT_465_data = 2'h0;
  assign mem_MPORT_465_addr = 9'h1d1;
  assign mem_MPORT_465_mask = 1'h1;
  assign mem_MPORT_465_en = reset;
  assign mem_MPORT_466_data = 2'h0;
  assign mem_MPORT_466_addr = 9'h1d2;
  assign mem_MPORT_466_mask = 1'h1;
  assign mem_MPORT_466_en = reset;
  assign mem_MPORT_467_data = 2'h0;
  assign mem_MPORT_467_addr = 9'h1d3;
  assign mem_MPORT_467_mask = 1'h1;
  assign mem_MPORT_467_en = reset;
  assign mem_MPORT_468_data = 2'h0;
  assign mem_MPORT_468_addr = 9'h1d4;
  assign mem_MPORT_468_mask = 1'h1;
  assign mem_MPORT_468_en = reset;
  assign mem_MPORT_469_data = 2'h0;
  assign mem_MPORT_469_addr = 9'h1d5;
  assign mem_MPORT_469_mask = 1'h1;
  assign mem_MPORT_469_en = reset;
  assign mem_MPORT_470_data = 2'h0;
  assign mem_MPORT_470_addr = 9'h1d6;
  assign mem_MPORT_470_mask = 1'h1;
  assign mem_MPORT_470_en = reset;
  assign mem_MPORT_471_data = 2'h0;
  assign mem_MPORT_471_addr = 9'h1d7;
  assign mem_MPORT_471_mask = 1'h1;
  assign mem_MPORT_471_en = reset;
  assign mem_MPORT_472_data = 2'h0;
  assign mem_MPORT_472_addr = 9'h1d8;
  assign mem_MPORT_472_mask = 1'h1;
  assign mem_MPORT_472_en = reset;
  assign mem_MPORT_473_data = 2'h0;
  assign mem_MPORT_473_addr = 9'h1d9;
  assign mem_MPORT_473_mask = 1'h1;
  assign mem_MPORT_473_en = reset;
  assign mem_MPORT_474_data = 2'h0;
  assign mem_MPORT_474_addr = 9'h1da;
  assign mem_MPORT_474_mask = 1'h1;
  assign mem_MPORT_474_en = reset;
  assign mem_MPORT_475_data = 2'h0;
  assign mem_MPORT_475_addr = 9'h1db;
  assign mem_MPORT_475_mask = 1'h1;
  assign mem_MPORT_475_en = reset;
  assign mem_MPORT_476_data = 2'h0;
  assign mem_MPORT_476_addr = 9'h1dc;
  assign mem_MPORT_476_mask = 1'h1;
  assign mem_MPORT_476_en = reset;
  assign mem_MPORT_477_data = 2'h0;
  assign mem_MPORT_477_addr = 9'h1dd;
  assign mem_MPORT_477_mask = 1'h1;
  assign mem_MPORT_477_en = reset;
  assign mem_MPORT_478_data = 2'h0;
  assign mem_MPORT_478_addr = 9'h1de;
  assign mem_MPORT_478_mask = 1'h1;
  assign mem_MPORT_478_en = reset;
  assign mem_MPORT_479_data = 2'h0;
  assign mem_MPORT_479_addr = 9'h1df;
  assign mem_MPORT_479_mask = 1'h1;
  assign mem_MPORT_479_en = reset;
  assign mem_MPORT_480_data = 2'h0;
  assign mem_MPORT_480_addr = 9'h1e0;
  assign mem_MPORT_480_mask = 1'h1;
  assign mem_MPORT_480_en = reset;
  assign mem_MPORT_481_data = 2'h0;
  assign mem_MPORT_481_addr = 9'h1e1;
  assign mem_MPORT_481_mask = 1'h1;
  assign mem_MPORT_481_en = reset;
  assign mem_MPORT_482_data = 2'h0;
  assign mem_MPORT_482_addr = 9'h1e2;
  assign mem_MPORT_482_mask = 1'h1;
  assign mem_MPORT_482_en = reset;
  assign mem_MPORT_483_data = 2'h0;
  assign mem_MPORT_483_addr = 9'h1e3;
  assign mem_MPORT_483_mask = 1'h1;
  assign mem_MPORT_483_en = reset;
  assign mem_MPORT_484_data = 2'h0;
  assign mem_MPORT_484_addr = 9'h1e4;
  assign mem_MPORT_484_mask = 1'h1;
  assign mem_MPORT_484_en = reset;
  assign mem_MPORT_485_data = 2'h0;
  assign mem_MPORT_485_addr = 9'h1e5;
  assign mem_MPORT_485_mask = 1'h1;
  assign mem_MPORT_485_en = reset;
  assign mem_MPORT_486_data = 2'h0;
  assign mem_MPORT_486_addr = 9'h1e6;
  assign mem_MPORT_486_mask = 1'h1;
  assign mem_MPORT_486_en = reset;
  assign mem_MPORT_487_data = 2'h0;
  assign mem_MPORT_487_addr = 9'h1e7;
  assign mem_MPORT_487_mask = 1'h1;
  assign mem_MPORT_487_en = reset;
  assign mem_MPORT_488_data = 2'h0;
  assign mem_MPORT_488_addr = 9'h1e8;
  assign mem_MPORT_488_mask = 1'h1;
  assign mem_MPORT_488_en = reset;
  assign mem_MPORT_489_data = 2'h0;
  assign mem_MPORT_489_addr = 9'h1e9;
  assign mem_MPORT_489_mask = 1'h1;
  assign mem_MPORT_489_en = reset;
  assign mem_MPORT_490_data = 2'h0;
  assign mem_MPORT_490_addr = 9'h1ea;
  assign mem_MPORT_490_mask = 1'h1;
  assign mem_MPORT_490_en = reset;
  assign mem_MPORT_491_data = 2'h0;
  assign mem_MPORT_491_addr = 9'h1eb;
  assign mem_MPORT_491_mask = 1'h1;
  assign mem_MPORT_491_en = reset;
  assign mem_MPORT_492_data = 2'h0;
  assign mem_MPORT_492_addr = 9'h1ec;
  assign mem_MPORT_492_mask = 1'h1;
  assign mem_MPORT_492_en = reset;
  assign mem_MPORT_493_data = 2'h0;
  assign mem_MPORT_493_addr = 9'h1ed;
  assign mem_MPORT_493_mask = 1'h1;
  assign mem_MPORT_493_en = reset;
  assign mem_MPORT_494_data = 2'h0;
  assign mem_MPORT_494_addr = 9'h1ee;
  assign mem_MPORT_494_mask = 1'h1;
  assign mem_MPORT_494_en = reset;
  assign mem_MPORT_495_data = 2'h0;
  assign mem_MPORT_495_addr = 9'h1ef;
  assign mem_MPORT_495_mask = 1'h1;
  assign mem_MPORT_495_en = reset;
  assign mem_MPORT_496_data = 2'h0;
  assign mem_MPORT_496_addr = 9'h1f0;
  assign mem_MPORT_496_mask = 1'h1;
  assign mem_MPORT_496_en = reset;
  assign mem_MPORT_497_data = 2'h0;
  assign mem_MPORT_497_addr = 9'h1f1;
  assign mem_MPORT_497_mask = 1'h1;
  assign mem_MPORT_497_en = reset;
  assign mem_MPORT_498_data = 2'h0;
  assign mem_MPORT_498_addr = 9'h1f2;
  assign mem_MPORT_498_mask = 1'h1;
  assign mem_MPORT_498_en = reset;
  assign mem_MPORT_499_data = 2'h0;
  assign mem_MPORT_499_addr = 9'h1f3;
  assign mem_MPORT_499_mask = 1'h1;
  assign mem_MPORT_499_en = reset;
  assign mem_MPORT_500_data = 2'h0;
  assign mem_MPORT_500_addr = 9'h1f4;
  assign mem_MPORT_500_mask = 1'h1;
  assign mem_MPORT_500_en = reset;
  assign mem_MPORT_501_data = 2'h0;
  assign mem_MPORT_501_addr = 9'h1f5;
  assign mem_MPORT_501_mask = 1'h1;
  assign mem_MPORT_501_en = reset;
  assign mem_MPORT_502_data = 2'h0;
  assign mem_MPORT_502_addr = 9'h1f6;
  assign mem_MPORT_502_mask = 1'h1;
  assign mem_MPORT_502_en = reset;
  assign mem_MPORT_503_data = 2'h0;
  assign mem_MPORT_503_addr = 9'h1f7;
  assign mem_MPORT_503_mask = 1'h1;
  assign mem_MPORT_503_en = reset;
  assign mem_MPORT_504_data = 2'h0;
  assign mem_MPORT_504_addr = 9'h1f8;
  assign mem_MPORT_504_mask = 1'h1;
  assign mem_MPORT_504_en = reset;
  assign mem_MPORT_505_data = 2'h0;
  assign mem_MPORT_505_addr = 9'h1f9;
  assign mem_MPORT_505_mask = 1'h1;
  assign mem_MPORT_505_en = reset;
  assign mem_MPORT_506_data = 2'h0;
  assign mem_MPORT_506_addr = 9'h1fa;
  assign mem_MPORT_506_mask = 1'h1;
  assign mem_MPORT_506_en = reset;
  assign mem_MPORT_507_data = 2'h0;
  assign mem_MPORT_507_addr = 9'h1fb;
  assign mem_MPORT_507_mask = 1'h1;
  assign mem_MPORT_507_en = reset;
  assign mem_MPORT_508_data = 2'h0;
  assign mem_MPORT_508_addr = 9'h1fc;
  assign mem_MPORT_508_mask = 1'h1;
  assign mem_MPORT_508_en = reset;
  assign mem_MPORT_509_data = 2'h0;
  assign mem_MPORT_509_addr = 9'h1fd;
  assign mem_MPORT_509_mask = 1'h1;
  assign mem_MPORT_509_en = reset;
  assign mem_MPORT_510_data = 2'h0;
  assign mem_MPORT_510_addr = 9'h1fe;
  assign mem_MPORT_510_mask = 1'h1;
  assign mem_MPORT_510_en = reset;
  assign mem_MPORT_511_data = 2'h0;
  assign mem_MPORT_511_addr = 9'h1ff;
  assign mem_MPORT_511_mask = 1'h1;
  assign mem_MPORT_511_en = reset;
  assign mem_MPORT_512_data = io_w_data;
  assign mem_MPORT_512_addr = io_w_addr;
  assign mem_MPORT_512_mask = 1'h1;
  assign mem_MPORT_512_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_129_en & mem_MPORT_129_mask) begin
      mem[mem_MPORT_129_addr] <= mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_130_en & mem_MPORT_130_mask) begin
      mem[mem_MPORT_130_addr] <= mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_131_en & mem_MPORT_131_mask) begin
      mem[mem_MPORT_131_addr] <= mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_132_en & mem_MPORT_132_mask) begin
      mem[mem_MPORT_132_addr] <= mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_133_en & mem_MPORT_133_mask) begin
      mem[mem_MPORT_133_addr] <= mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_134_en & mem_MPORT_134_mask) begin
      mem[mem_MPORT_134_addr] <= mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_135_en & mem_MPORT_135_mask) begin
      mem[mem_MPORT_135_addr] <= mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_136_en & mem_MPORT_136_mask) begin
      mem[mem_MPORT_136_addr] <= mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_137_en & mem_MPORT_137_mask) begin
      mem[mem_MPORT_137_addr] <= mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_138_en & mem_MPORT_138_mask) begin
      mem[mem_MPORT_138_addr] <= mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_139_en & mem_MPORT_139_mask) begin
      mem[mem_MPORT_139_addr] <= mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_140_en & mem_MPORT_140_mask) begin
      mem[mem_MPORT_140_addr] <= mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_141_en & mem_MPORT_141_mask) begin
      mem[mem_MPORT_141_addr] <= mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_142_en & mem_MPORT_142_mask) begin
      mem[mem_MPORT_142_addr] <= mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_143_en & mem_MPORT_143_mask) begin
      mem[mem_MPORT_143_addr] <= mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_144_en & mem_MPORT_144_mask) begin
      mem[mem_MPORT_144_addr] <= mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_145_en & mem_MPORT_145_mask) begin
      mem[mem_MPORT_145_addr] <= mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_146_en & mem_MPORT_146_mask) begin
      mem[mem_MPORT_146_addr] <= mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_147_en & mem_MPORT_147_mask) begin
      mem[mem_MPORT_147_addr] <= mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_148_en & mem_MPORT_148_mask) begin
      mem[mem_MPORT_148_addr] <= mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_149_en & mem_MPORT_149_mask) begin
      mem[mem_MPORT_149_addr] <= mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_150_en & mem_MPORT_150_mask) begin
      mem[mem_MPORT_150_addr] <= mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_151_en & mem_MPORT_151_mask) begin
      mem[mem_MPORT_151_addr] <= mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_152_en & mem_MPORT_152_mask) begin
      mem[mem_MPORT_152_addr] <= mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_153_en & mem_MPORT_153_mask) begin
      mem[mem_MPORT_153_addr] <= mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_154_en & mem_MPORT_154_mask) begin
      mem[mem_MPORT_154_addr] <= mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_155_en & mem_MPORT_155_mask) begin
      mem[mem_MPORT_155_addr] <= mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_156_en & mem_MPORT_156_mask) begin
      mem[mem_MPORT_156_addr] <= mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_157_en & mem_MPORT_157_mask) begin
      mem[mem_MPORT_157_addr] <= mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_158_en & mem_MPORT_158_mask) begin
      mem[mem_MPORT_158_addr] <= mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_159_en & mem_MPORT_159_mask) begin
      mem[mem_MPORT_159_addr] <= mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_160_en & mem_MPORT_160_mask) begin
      mem[mem_MPORT_160_addr] <= mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_161_en & mem_MPORT_161_mask) begin
      mem[mem_MPORT_161_addr] <= mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_162_en & mem_MPORT_162_mask) begin
      mem[mem_MPORT_162_addr] <= mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_163_en & mem_MPORT_163_mask) begin
      mem[mem_MPORT_163_addr] <= mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_164_en & mem_MPORT_164_mask) begin
      mem[mem_MPORT_164_addr] <= mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_165_en & mem_MPORT_165_mask) begin
      mem[mem_MPORT_165_addr] <= mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_166_en & mem_MPORT_166_mask) begin
      mem[mem_MPORT_166_addr] <= mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_167_en & mem_MPORT_167_mask) begin
      mem[mem_MPORT_167_addr] <= mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_168_en & mem_MPORT_168_mask) begin
      mem[mem_MPORT_168_addr] <= mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_169_en & mem_MPORT_169_mask) begin
      mem[mem_MPORT_169_addr] <= mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_170_en & mem_MPORT_170_mask) begin
      mem[mem_MPORT_170_addr] <= mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_171_en & mem_MPORT_171_mask) begin
      mem[mem_MPORT_171_addr] <= mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_172_en & mem_MPORT_172_mask) begin
      mem[mem_MPORT_172_addr] <= mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_173_en & mem_MPORT_173_mask) begin
      mem[mem_MPORT_173_addr] <= mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_174_en & mem_MPORT_174_mask) begin
      mem[mem_MPORT_174_addr] <= mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_175_en & mem_MPORT_175_mask) begin
      mem[mem_MPORT_175_addr] <= mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_176_en & mem_MPORT_176_mask) begin
      mem[mem_MPORT_176_addr] <= mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_177_en & mem_MPORT_177_mask) begin
      mem[mem_MPORT_177_addr] <= mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_178_en & mem_MPORT_178_mask) begin
      mem[mem_MPORT_178_addr] <= mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_179_en & mem_MPORT_179_mask) begin
      mem[mem_MPORT_179_addr] <= mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_180_en & mem_MPORT_180_mask) begin
      mem[mem_MPORT_180_addr] <= mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_181_en & mem_MPORT_181_mask) begin
      mem[mem_MPORT_181_addr] <= mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_182_en & mem_MPORT_182_mask) begin
      mem[mem_MPORT_182_addr] <= mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_183_en & mem_MPORT_183_mask) begin
      mem[mem_MPORT_183_addr] <= mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_184_en & mem_MPORT_184_mask) begin
      mem[mem_MPORT_184_addr] <= mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_185_en & mem_MPORT_185_mask) begin
      mem[mem_MPORT_185_addr] <= mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_186_en & mem_MPORT_186_mask) begin
      mem[mem_MPORT_186_addr] <= mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_187_en & mem_MPORT_187_mask) begin
      mem[mem_MPORT_187_addr] <= mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_188_en & mem_MPORT_188_mask) begin
      mem[mem_MPORT_188_addr] <= mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_189_en & mem_MPORT_189_mask) begin
      mem[mem_MPORT_189_addr] <= mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_190_en & mem_MPORT_190_mask) begin
      mem[mem_MPORT_190_addr] <= mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_191_en & mem_MPORT_191_mask) begin
      mem[mem_MPORT_191_addr] <= mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_192_en & mem_MPORT_192_mask) begin
      mem[mem_MPORT_192_addr] <= mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_193_en & mem_MPORT_193_mask) begin
      mem[mem_MPORT_193_addr] <= mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_194_en & mem_MPORT_194_mask) begin
      mem[mem_MPORT_194_addr] <= mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_195_en & mem_MPORT_195_mask) begin
      mem[mem_MPORT_195_addr] <= mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_196_en & mem_MPORT_196_mask) begin
      mem[mem_MPORT_196_addr] <= mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_197_en & mem_MPORT_197_mask) begin
      mem[mem_MPORT_197_addr] <= mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_198_en & mem_MPORT_198_mask) begin
      mem[mem_MPORT_198_addr] <= mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_199_en & mem_MPORT_199_mask) begin
      mem[mem_MPORT_199_addr] <= mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_200_en & mem_MPORT_200_mask) begin
      mem[mem_MPORT_200_addr] <= mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_201_en & mem_MPORT_201_mask) begin
      mem[mem_MPORT_201_addr] <= mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_202_en & mem_MPORT_202_mask) begin
      mem[mem_MPORT_202_addr] <= mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_203_en & mem_MPORT_203_mask) begin
      mem[mem_MPORT_203_addr] <= mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_204_en & mem_MPORT_204_mask) begin
      mem[mem_MPORT_204_addr] <= mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_205_en & mem_MPORT_205_mask) begin
      mem[mem_MPORT_205_addr] <= mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_206_en & mem_MPORT_206_mask) begin
      mem[mem_MPORT_206_addr] <= mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_207_en & mem_MPORT_207_mask) begin
      mem[mem_MPORT_207_addr] <= mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_208_en & mem_MPORT_208_mask) begin
      mem[mem_MPORT_208_addr] <= mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_209_en & mem_MPORT_209_mask) begin
      mem[mem_MPORT_209_addr] <= mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_210_en & mem_MPORT_210_mask) begin
      mem[mem_MPORT_210_addr] <= mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_211_en & mem_MPORT_211_mask) begin
      mem[mem_MPORT_211_addr] <= mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_212_en & mem_MPORT_212_mask) begin
      mem[mem_MPORT_212_addr] <= mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_213_en & mem_MPORT_213_mask) begin
      mem[mem_MPORT_213_addr] <= mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_214_en & mem_MPORT_214_mask) begin
      mem[mem_MPORT_214_addr] <= mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_215_en & mem_MPORT_215_mask) begin
      mem[mem_MPORT_215_addr] <= mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_216_en & mem_MPORT_216_mask) begin
      mem[mem_MPORT_216_addr] <= mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_217_en & mem_MPORT_217_mask) begin
      mem[mem_MPORT_217_addr] <= mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_218_en & mem_MPORT_218_mask) begin
      mem[mem_MPORT_218_addr] <= mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_219_en & mem_MPORT_219_mask) begin
      mem[mem_MPORT_219_addr] <= mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_220_en & mem_MPORT_220_mask) begin
      mem[mem_MPORT_220_addr] <= mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_221_en & mem_MPORT_221_mask) begin
      mem[mem_MPORT_221_addr] <= mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_222_en & mem_MPORT_222_mask) begin
      mem[mem_MPORT_222_addr] <= mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_223_en & mem_MPORT_223_mask) begin
      mem[mem_MPORT_223_addr] <= mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_224_en & mem_MPORT_224_mask) begin
      mem[mem_MPORT_224_addr] <= mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_225_en & mem_MPORT_225_mask) begin
      mem[mem_MPORT_225_addr] <= mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_226_en & mem_MPORT_226_mask) begin
      mem[mem_MPORT_226_addr] <= mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_227_en & mem_MPORT_227_mask) begin
      mem[mem_MPORT_227_addr] <= mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_228_en & mem_MPORT_228_mask) begin
      mem[mem_MPORT_228_addr] <= mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_229_en & mem_MPORT_229_mask) begin
      mem[mem_MPORT_229_addr] <= mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_230_en & mem_MPORT_230_mask) begin
      mem[mem_MPORT_230_addr] <= mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_231_en & mem_MPORT_231_mask) begin
      mem[mem_MPORT_231_addr] <= mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_232_en & mem_MPORT_232_mask) begin
      mem[mem_MPORT_232_addr] <= mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_233_en & mem_MPORT_233_mask) begin
      mem[mem_MPORT_233_addr] <= mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_234_en & mem_MPORT_234_mask) begin
      mem[mem_MPORT_234_addr] <= mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_235_en & mem_MPORT_235_mask) begin
      mem[mem_MPORT_235_addr] <= mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_236_en & mem_MPORT_236_mask) begin
      mem[mem_MPORT_236_addr] <= mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_237_en & mem_MPORT_237_mask) begin
      mem[mem_MPORT_237_addr] <= mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_238_en & mem_MPORT_238_mask) begin
      mem[mem_MPORT_238_addr] <= mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_239_en & mem_MPORT_239_mask) begin
      mem[mem_MPORT_239_addr] <= mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_240_en & mem_MPORT_240_mask) begin
      mem[mem_MPORT_240_addr] <= mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_241_en & mem_MPORT_241_mask) begin
      mem[mem_MPORT_241_addr] <= mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_242_en & mem_MPORT_242_mask) begin
      mem[mem_MPORT_242_addr] <= mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_243_en & mem_MPORT_243_mask) begin
      mem[mem_MPORT_243_addr] <= mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_244_en & mem_MPORT_244_mask) begin
      mem[mem_MPORT_244_addr] <= mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_245_en & mem_MPORT_245_mask) begin
      mem[mem_MPORT_245_addr] <= mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_246_en & mem_MPORT_246_mask) begin
      mem[mem_MPORT_246_addr] <= mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_247_en & mem_MPORT_247_mask) begin
      mem[mem_MPORT_247_addr] <= mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_248_en & mem_MPORT_248_mask) begin
      mem[mem_MPORT_248_addr] <= mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_249_en & mem_MPORT_249_mask) begin
      mem[mem_MPORT_249_addr] <= mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_250_en & mem_MPORT_250_mask) begin
      mem[mem_MPORT_250_addr] <= mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_251_en & mem_MPORT_251_mask) begin
      mem[mem_MPORT_251_addr] <= mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_252_en & mem_MPORT_252_mask) begin
      mem[mem_MPORT_252_addr] <= mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_253_en & mem_MPORT_253_mask) begin
      mem[mem_MPORT_253_addr] <= mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_254_en & mem_MPORT_254_mask) begin
      mem[mem_MPORT_254_addr] <= mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_255_en & mem_MPORT_255_mask) begin
      mem[mem_MPORT_255_addr] <= mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_256_en & mem_MPORT_256_mask) begin
      mem[mem_MPORT_256_addr] <= mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_257_en & mem_MPORT_257_mask) begin
      mem[mem_MPORT_257_addr] <= mem_MPORT_257_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_258_en & mem_MPORT_258_mask) begin
      mem[mem_MPORT_258_addr] <= mem_MPORT_258_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_259_en & mem_MPORT_259_mask) begin
      mem[mem_MPORT_259_addr] <= mem_MPORT_259_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_260_en & mem_MPORT_260_mask) begin
      mem[mem_MPORT_260_addr] <= mem_MPORT_260_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_261_en & mem_MPORT_261_mask) begin
      mem[mem_MPORT_261_addr] <= mem_MPORT_261_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_262_en & mem_MPORT_262_mask) begin
      mem[mem_MPORT_262_addr] <= mem_MPORT_262_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_263_en & mem_MPORT_263_mask) begin
      mem[mem_MPORT_263_addr] <= mem_MPORT_263_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_264_en & mem_MPORT_264_mask) begin
      mem[mem_MPORT_264_addr] <= mem_MPORT_264_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_265_en & mem_MPORT_265_mask) begin
      mem[mem_MPORT_265_addr] <= mem_MPORT_265_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_266_en & mem_MPORT_266_mask) begin
      mem[mem_MPORT_266_addr] <= mem_MPORT_266_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_267_en & mem_MPORT_267_mask) begin
      mem[mem_MPORT_267_addr] <= mem_MPORT_267_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_268_en & mem_MPORT_268_mask) begin
      mem[mem_MPORT_268_addr] <= mem_MPORT_268_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_269_en & mem_MPORT_269_mask) begin
      mem[mem_MPORT_269_addr] <= mem_MPORT_269_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_270_en & mem_MPORT_270_mask) begin
      mem[mem_MPORT_270_addr] <= mem_MPORT_270_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_271_en & mem_MPORT_271_mask) begin
      mem[mem_MPORT_271_addr] <= mem_MPORT_271_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_272_en & mem_MPORT_272_mask) begin
      mem[mem_MPORT_272_addr] <= mem_MPORT_272_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_273_en & mem_MPORT_273_mask) begin
      mem[mem_MPORT_273_addr] <= mem_MPORT_273_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_274_en & mem_MPORT_274_mask) begin
      mem[mem_MPORT_274_addr] <= mem_MPORT_274_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_275_en & mem_MPORT_275_mask) begin
      mem[mem_MPORT_275_addr] <= mem_MPORT_275_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_276_en & mem_MPORT_276_mask) begin
      mem[mem_MPORT_276_addr] <= mem_MPORT_276_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_277_en & mem_MPORT_277_mask) begin
      mem[mem_MPORT_277_addr] <= mem_MPORT_277_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_278_en & mem_MPORT_278_mask) begin
      mem[mem_MPORT_278_addr] <= mem_MPORT_278_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_279_en & mem_MPORT_279_mask) begin
      mem[mem_MPORT_279_addr] <= mem_MPORT_279_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_280_en & mem_MPORT_280_mask) begin
      mem[mem_MPORT_280_addr] <= mem_MPORT_280_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_281_en & mem_MPORT_281_mask) begin
      mem[mem_MPORT_281_addr] <= mem_MPORT_281_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_282_en & mem_MPORT_282_mask) begin
      mem[mem_MPORT_282_addr] <= mem_MPORT_282_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_283_en & mem_MPORT_283_mask) begin
      mem[mem_MPORT_283_addr] <= mem_MPORT_283_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_284_en & mem_MPORT_284_mask) begin
      mem[mem_MPORT_284_addr] <= mem_MPORT_284_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_285_en & mem_MPORT_285_mask) begin
      mem[mem_MPORT_285_addr] <= mem_MPORT_285_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_286_en & mem_MPORT_286_mask) begin
      mem[mem_MPORT_286_addr] <= mem_MPORT_286_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_287_en & mem_MPORT_287_mask) begin
      mem[mem_MPORT_287_addr] <= mem_MPORT_287_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_288_en & mem_MPORT_288_mask) begin
      mem[mem_MPORT_288_addr] <= mem_MPORT_288_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_289_en & mem_MPORT_289_mask) begin
      mem[mem_MPORT_289_addr] <= mem_MPORT_289_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_290_en & mem_MPORT_290_mask) begin
      mem[mem_MPORT_290_addr] <= mem_MPORT_290_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_291_en & mem_MPORT_291_mask) begin
      mem[mem_MPORT_291_addr] <= mem_MPORT_291_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_292_en & mem_MPORT_292_mask) begin
      mem[mem_MPORT_292_addr] <= mem_MPORT_292_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_293_en & mem_MPORT_293_mask) begin
      mem[mem_MPORT_293_addr] <= mem_MPORT_293_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_294_en & mem_MPORT_294_mask) begin
      mem[mem_MPORT_294_addr] <= mem_MPORT_294_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_295_en & mem_MPORT_295_mask) begin
      mem[mem_MPORT_295_addr] <= mem_MPORT_295_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_296_en & mem_MPORT_296_mask) begin
      mem[mem_MPORT_296_addr] <= mem_MPORT_296_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_297_en & mem_MPORT_297_mask) begin
      mem[mem_MPORT_297_addr] <= mem_MPORT_297_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_298_en & mem_MPORT_298_mask) begin
      mem[mem_MPORT_298_addr] <= mem_MPORT_298_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_299_en & mem_MPORT_299_mask) begin
      mem[mem_MPORT_299_addr] <= mem_MPORT_299_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_300_en & mem_MPORT_300_mask) begin
      mem[mem_MPORT_300_addr] <= mem_MPORT_300_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_301_en & mem_MPORT_301_mask) begin
      mem[mem_MPORT_301_addr] <= mem_MPORT_301_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_302_en & mem_MPORT_302_mask) begin
      mem[mem_MPORT_302_addr] <= mem_MPORT_302_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_303_en & mem_MPORT_303_mask) begin
      mem[mem_MPORT_303_addr] <= mem_MPORT_303_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_304_en & mem_MPORT_304_mask) begin
      mem[mem_MPORT_304_addr] <= mem_MPORT_304_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_305_en & mem_MPORT_305_mask) begin
      mem[mem_MPORT_305_addr] <= mem_MPORT_305_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_306_en & mem_MPORT_306_mask) begin
      mem[mem_MPORT_306_addr] <= mem_MPORT_306_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_307_en & mem_MPORT_307_mask) begin
      mem[mem_MPORT_307_addr] <= mem_MPORT_307_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_308_en & mem_MPORT_308_mask) begin
      mem[mem_MPORT_308_addr] <= mem_MPORT_308_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_309_en & mem_MPORT_309_mask) begin
      mem[mem_MPORT_309_addr] <= mem_MPORT_309_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_310_en & mem_MPORT_310_mask) begin
      mem[mem_MPORT_310_addr] <= mem_MPORT_310_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_311_en & mem_MPORT_311_mask) begin
      mem[mem_MPORT_311_addr] <= mem_MPORT_311_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_312_en & mem_MPORT_312_mask) begin
      mem[mem_MPORT_312_addr] <= mem_MPORT_312_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_313_en & mem_MPORT_313_mask) begin
      mem[mem_MPORT_313_addr] <= mem_MPORT_313_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_314_en & mem_MPORT_314_mask) begin
      mem[mem_MPORT_314_addr] <= mem_MPORT_314_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_315_en & mem_MPORT_315_mask) begin
      mem[mem_MPORT_315_addr] <= mem_MPORT_315_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_316_en & mem_MPORT_316_mask) begin
      mem[mem_MPORT_316_addr] <= mem_MPORT_316_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_317_en & mem_MPORT_317_mask) begin
      mem[mem_MPORT_317_addr] <= mem_MPORT_317_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_318_en & mem_MPORT_318_mask) begin
      mem[mem_MPORT_318_addr] <= mem_MPORT_318_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_319_en & mem_MPORT_319_mask) begin
      mem[mem_MPORT_319_addr] <= mem_MPORT_319_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_320_en & mem_MPORT_320_mask) begin
      mem[mem_MPORT_320_addr] <= mem_MPORT_320_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_321_en & mem_MPORT_321_mask) begin
      mem[mem_MPORT_321_addr] <= mem_MPORT_321_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_322_en & mem_MPORT_322_mask) begin
      mem[mem_MPORT_322_addr] <= mem_MPORT_322_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_323_en & mem_MPORT_323_mask) begin
      mem[mem_MPORT_323_addr] <= mem_MPORT_323_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_324_en & mem_MPORT_324_mask) begin
      mem[mem_MPORT_324_addr] <= mem_MPORT_324_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_325_en & mem_MPORT_325_mask) begin
      mem[mem_MPORT_325_addr] <= mem_MPORT_325_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_326_en & mem_MPORT_326_mask) begin
      mem[mem_MPORT_326_addr] <= mem_MPORT_326_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_327_en & mem_MPORT_327_mask) begin
      mem[mem_MPORT_327_addr] <= mem_MPORT_327_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_328_en & mem_MPORT_328_mask) begin
      mem[mem_MPORT_328_addr] <= mem_MPORT_328_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_329_en & mem_MPORT_329_mask) begin
      mem[mem_MPORT_329_addr] <= mem_MPORT_329_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_330_en & mem_MPORT_330_mask) begin
      mem[mem_MPORT_330_addr] <= mem_MPORT_330_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_331_en & mem_MPORT_331_mask) begin
      mem[mem_MPORT_331_addr] <= mem_MPORT_331_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_332_en & mem_MPORT_332_mask) begin
      mem[mem_MPORT_332_addr] <= mem_MPORT_332_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_333_en & mem_MPORT_333_mask) begin
      mem[mem_MPORT_333_addr] <= mem_MPORT_333_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_334_en & mem_MPORT_334_mask) begin
      mem[mem_MPORT_334_addr] <= mem_MPORT_334_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_335_en & mem_MPORT_335_mask) begin
      mem[mem_MPORT_335_addr] <= mem_MPORT_335_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_336_en & mem_MPORT_336_mask) begin
      mem[mem_MPORT_336_addr] <= mem_MPORT_336_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_337_en & mem_MPORT_337_mask) begin
      mem[mem_MPORT_337_addr] <= mem_MPORT_337_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_338_en & mem_MPORT_338_mask) begin
      mem[mem_MPORT_338_addr] <= mem_MPORT_338_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_339_en & mem_MPORT_339_mask) begin
      mem[mem_MPORT_339_addr] <= mem_MPORT_339_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_340_en & mem_MPORT_340_mask) begin
      mem[mem_MPORT_340_addr] <= mem_MPORT_340_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_341_en & mem_MPORT_341_mask) begin
      mem[mem_MPORT_341_addr] <= mem_MPORT_341_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_342_en & mem_MPORT_342_mask) begin
      mem[mem_MPORT_342_addr] <= mem_MPORT_342_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_343_en & mem_MPORT_343_mask) begin
      mem[mem_MPORT_343_addr] <= mem_MPORT_343_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_344_en & mem_MPORT_344_mask) begin
      mem[mem_MPORT_344_addr] <= mem_MPORT_344_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_345_en & mem_MPORT_345_mask) begin
      mem[mem_MPORT_345_addr] <= mem_MPORT_345_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_346_en & mem_MPORT_346_mask) begin
      mem[mem_MPORT_346_addr] <= mem_MPORT_346_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_347_en & mem_MPORT_347_mask) begin
      mem[mem_MPORT_347_addr] <= mem_MPORT_347_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_348_en & mem_MPORT_348_mask) begin
      mem[mem_MPORT_348_addr] <= mem_MPORT_348_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_349_en & mem_MPORT_349_mask) begin
      mem[mem_MPORT_349_addr] <= mem_MPORT_349_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_350_en & mem_MPORT_350_mask) begin
      mem[mem_MPORT_350_addr] <= mem_MPORT_350_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_351_en & mem_MPORT_351_mask) begin
      mem[mem_MPORT_351_addr] <= mem_MPORT_351_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_352_en & mem_MPORT_352_mask) begin
      mem[mem_MPORT_352_addr] <= mem_MPORT_352_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_353_en & mem_MPORT_353_mask) begin
      mem[mem_MPORT_353_addr] <= mem_MPORT_353_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_354_en & mem_MPORT_354_mask) begin
      mem[mem_MPORT_354_addr] <= mem_MPORT_354_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_355_en & mem_MPORT_355_mask) begin
      mem[mem_MPORT_355_addr] <= mem_MPORT_355_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_356_en & mem_MPORT_356_mask) begin
      mem[mem_MPORT_356_addr] <= mem_MPORT_356_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_357_en & mem_MPORT_357_mask) begin
      mem[mem_MPORT_357_addr] <= mem_MPORT_357_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_358_en & mem_MPORT_358_mask) begin
      mem[mem_MPORT_358_addr] <= mem_MPORT_358_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_359_en & mem_MPORT_359_mask) begin
      mem[mem_MPORT_359_addr] <= mem_MPORT_359_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_360_en & mem_MPORT_360_mask) begin
      mem[mem_MPORT_360_addr] <= mem_MPORT_360_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_361_en & mem_MPORT_361_mask) begin
      mem[mem_MPORT_361_addr] <= mem_MPORT_361_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_362_en & mem_MPORT_362_mask) begin
      mem[mem_MPORT_362_addr] <= mem_MPORT_362_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_363_en & mem_MPORT_363_mask) begin
      mem[mem_MPORT_363_addr] <= mem_MPORT_363_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_364_en & mem_MPORT_364_mask) begin
      mem[mem_MPORT_364_addr] <= mem_MPORT_364_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_365_en & mem_MPORT_365_mask) begin
      mem[mem_MPORT_365_addr] <= mem_MPORT_365_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_366_en & mem_MPORT_366_mask) begin
      mem[mem_MPORT_366_addr] <= mem_MPORT_366_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_367_en & mem_MPORT_367_mask) begin
      mem[mem_MPORT_367_addr] <= mem_MPORT_367_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_368_en & mem_MPORT_368_mask) begin
      mem[mem_MPORT_368_addr] <= mem_MPORT_368_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_369_en & mem_MPORT_369_mask) begin
      mem[mem_MPORT_369_addr] <= mem_MPORT_369_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_370_en & mem_MPORT_370_mask) begin
      mem[mem_MPORT_370_addr] <= mem_MPORT_370_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_371_en & mem_MPORT_371_mask) begin
      mem[mem_MPORT_371_addr] <= mem_MPORT_371_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_372_en & mem_MPORT_372_mask) begin
      mem[mem_MPORT_372_addr] <= mem_MPORT_372_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_373_en & mem_MPORT_373_mask) begin
      mem[mem_MPORT_373_addr] <= mem_MPORT_373_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_374_en & mem_MPORT_374_mask) begin
      mem[mem_MPORT_374_addr] <= mem_MPORT_374_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_375_en & mem_MPORT_375_mask) begin
      mem[mem_MPORT_375_addr] <= mem_MPORT_375_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_376_en & mem_MPORT_376_mask) begin
      mem[mem_MPORT_376_addr] <= mem_MPORT_376_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_377_en & mem_MPORT_377_mask) begin
      mem[mem_MPORT_377_addr] <= mem_MPORT_377_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_378_en & mem_MPORT_378_mask) begin
      mem[mem_MPORT_378_addr] <= mem_MPORT_378_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_379_en & mem_MPORT_379_mask) begin
      mem[mem_MPORT_379_addr] <= mem_MPORT_379_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_380_en & mem_MPORT_380_mask) begin
      mem[mem_MPORT_380_addr] <= mem_MPORT_380_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_381_en & mem_MPORT_381_mask) begin
      mem[mem_MPORT_381_addr] <= mem_MPORT_381_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_382_en & mem_MPORT_382_mask) begin
      mem[mem_MPORT_382_addr] <= mem_MPORT_382_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_383_en & mem_MPORT_383_mask) begin
      mem[mem_MPORT_383_addr] <= mem_MPORT_383_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_384_en & mem_MPORT_384_mask) begin
      mem[mem_MPORT_384_addr] <= mem_MPORT_384_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_385_en & mem_MPORT_385_mask) begin
      mem[mem_MPORT_385_addr] <= mem_MPORT_385_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_386_en & mem_MPORT_386_mask) begin
      mem[mem_MPORT_386_addr] <= mem_MPORT_386_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_387_en & mem_MPORT_387_mask) begin
      mem[mem_MPORT_387_addr] <= mem_MPORT_387_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_388_en & mem_MPORT_388_mask) begin
      mem[mem_MPORT_388_addr] <= mem_MPORT_388_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_389_en & mem_MPORT_389_mask) begin
      mem[mem_MPORT_389_addr] <= mem_MPORT_389_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_390_en & mem_MPORT_390_mask) begin
      mem[mem_MPORT_390_addr] <= mem_MPORT_390_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_391_en & mem_MPORT_391_mask) begin
      mem[mem_MPORT_391_addr] <= mem_MPORT_391_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_392_en & mem_MPORT_392_mask) begin
      mem[mem_MPORT_392_addr] <= mem_MPORT_392_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_393_en & mem_MPORT_393_mask) begin
      mem[mem_MPORT_393_addr] <= mem_MPORT_393_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_394_en & mem_MPORT_394_mask) begin
      mem[mem_MPORT_394_addr] <= mem_MPORT_394_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_395_en & mem_MPORT_395_mask) begin
      mem[mem_MPORT_395_addr] <= mem_MPORT_395_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_396_en & mem_MPORT_396_mask) begin
      mem[mem_MPORT_396_addr] <= mem_MPORT_396_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_397_en & mem_MPORT_397_mask) begin
      mem[mem_MPORT_397_addr] <= mem_MPORT_397_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_398_en & mem_MPORT_398_mask) begin
      mem[mem_MPORT_398_addr] <= mem_MPORT_398_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_399_en & mem_MPORT_399_mask) begin
      mem[mem_MPORT_399_addr] <= mem_MPORT_399_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_400_en & mem_MPORT_400_mask) begin
      mem[mem_MPORT_400_addr] <= mem_MPORT_400_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_401_en & mem_MPORT_401_mask) begin
      mem[mem_MPORT_401_addr] <= mem_MPORT_401_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_402_en & mem_MPORT_402_mask) begin
      mem[mem_MPORT_402_addr] <= mem_MPORT_402_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_403_en & mem_MPORT_403_mask) begin
      mem[mem_MPORT_403_addr] <= mem_MPORT_403_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_404_en & mem_MPORT_404_mask) begin
      mem[mem_MPORT_404_addr] <= mem_MPORT_404_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_405_en & mem_MPORT_405_mask) begin
      mem[mem_MPORT_405_addr] <= mem_MPORT_405_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_406_en & mem_MPORT_406_mask) begin
      mem[mem_MPORT_406_addr] <= mem_MPORT_406_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_407_en & mem_MPORT_407_mask) begin
      mem[mem_MPORT_407_addr] <= mem_MPORT_407_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_408_en & mem_MPORT_408_mask) begin
      mem[mem_MPORT_408_addr] <= mem_MPORT_408_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_409_en & mem_MPORT_409_mask) begin
      mem[mem_MPORT_409_addr] <= mem_MPORT_409_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_410_en & mem_MPORT_410_mask) begin
      mem[mem_MPORT_410_addr] <= mem_MPORT_410_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_411_en & mem_MPORT_411_mask) begin
      mem[mem_MPORT_411_addr] <= mem_MPORT_411_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_412_en & mem_MPORT_412_mask) begin
      mem[mem_MPORT_412_addr] <= mem_MPORT_412_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_413_en & mem_MPORT_413_mask) begin
      mem[mem_MPORT_413_addr] <= mem_MPORT_413_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_414_en & mem_MPORT_414_mask) begin
      mem[mem_MPORT_414_addr] <= mem_MPORT_414_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_415_en & mem_MPORT_415_mask) begin
      mem[mem_MPORT_415_addr] <= mem_MPORT_415_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_416_en & mem_MPORT_416_mask) begin
      mem[mem_MPORT_416_addr] <= mem_MPORT_416_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_417_en & mem_MPORT_417_mask) begin
      mem[mem_MPORT_417_addr] <= mem_MPORT_417_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_418_en & mem_MPORT_418_mask) begin
      mem[mem_MPORT_418_addr] <= mem_MPORT_418_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_419_en & mem_MPORT_419_mask) begin
      mem[mem_MPORT_419_addr] <= mem_MPORT_419_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_420_en & mem_MPORT_420_mask) begin
      mem[mem_MPORT_420_addr] <= mem_MPORT_420_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_421_en & mem_MPORT_421_mask) begin
      mem[mem_MPORT_421_addr] <= mem_MPORT_421_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_422_en & mem_MPORT_422_mask) begin
      mem[mem_MPORT_422_addr] <= mem_MPORT_422_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_423_en & mem_MPORT_423_mask) begin
      mem[mem_MPORT_423_addr] <= mem_MPORT_423_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_424_en & mem_MPORT_424_mask) begin
      mem[mem_MPORT_424_addr] <= mem_MPORT_424_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_425_en & mem_MPORT_425_mask) begin
      mem[mem_MPORT_425_addr] <= mem_MPORT_425_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_426_en & mem_MPORT_426_mask) begin
      mem[mem_MPORT_426_addr] <= mem_MPORT_426_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_427_en & mem_MPORT_427_mask) begin
      mem[mem_MPORT_427_addr] <= mem_MPORT_427_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_428_en & mem_MPORT_428_mask) begin
      mem[mem_MPORT_428_addr] <= mem_MPORT_428_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_429_en & mem_MPORT_429_mask) begin
      mem[mem_MPORT_429_addr] <= mem_MPORT_429_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_430_en & mem_MPORT_430_mask) begin
      mem[mem_MPORT_430_addr] <= mem_MPORT_430_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_431_en & mem_MPORT_431_mask) begin
      mem[mem_MPORT_431_addr] <= mem_MPORT_431_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_432_en & mem_MPORT_432_mask) begin
      mem[mem_MPORT_432_addr] <= mem_MPORT_432_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_433_en & mem_MPORT_433_mask) begin
      mem[mem_MPORT_433_addr] <= mem_MPORT_433_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_434_en & mem_MPORT_434_mask) begin
      mem[mem_MPORT_434_addr] <= mem_MPORT_434_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_435_en & mem_MPORT_435_mask) begin
      mem[mem_MPORT_435_addr] <= mem_MPORT_435_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_436_en & mem_MPORT_436_mask) begin
      mem[mem_MPORT_436_addr] <= mem_MPORT_436_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_437_en & mem_MPORT_437_mask) begin
      mem[mem_MPORT_437_addr] <= mem_MPORT_437_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_438_en & mem_MPORT_438_mask) begin
      mem[mem_MPORT_438_addr] <= mem_MPORT_438_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_439_en & mem_MPORT_439_mask) begin
      mem[mem_MPORT_439_addr] <= mem_MPORT_439_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_440_en & mem_MPORT_440_mask) begin
      mem[mem_MPORT_440_addr] <= mem_MPORT_440_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_441_en & mem_MPORT_441_mask) begin
      mem[mem_MPORT_441_addr] <= mem_MPORT_441_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_442_en & mem_MPORT_442_mask) begin
      mem[mem_MPORT_442_addr] <= mem_MPORT_442_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_443_en & mem_MPORT_443_mask) begin
      mem[mem_MPORT_443_addr] <= mem_MPORT_443_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_444_en & mem_MPORT_444_mask) begin
      mem[mem_MPORT_444_addr] <= mem_MPORT_444_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_445_en & mem_MPORT_445_mask) begin
      mem[mem_MPORT_445_addr] <= mem_MPORT_445_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_446_en & mem_MPORT_446_mask) begin
      mem[mem_MPORT_446_addr] <= mem_MPORT_446_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_447_en & mem_MPORT_447_mask) begin
      mem[mem_MPORT_447_addr] <= mem_MPORT_447_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_448_en & mem_MPORT_448_mask) begin
      mem[mem_MPORT_448_addr] <= mem_MPORT_448_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_449_en & mem_MPORT_449_mask) begin
      mem[mem_MPORT_449_addr] <= mem_MPORT_449_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_450_en & mem_MPORT_450_mask) begin
      mem[mem_MPORT_450_addr] <= mem_MPORT_450_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_451_en & mem_MPORT_451_mask) begin
      mem[mem_MPORT_451_addr] <= mem_MPORT_451_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_452_en & mem_MPORT_452_mask) begin
      mem[mem_MPORT_452_addr] <= mem_MPORT_452_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_453_en & mem_MPORT_453_mask) begin
      mem[mem_MPORT_453_addr] <= mem_MPORT_453_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_454_en & mem_MPORT_454_mask) begin
      mem[mem_MPORT_454_addr] <= mem_MPORT_454_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_455_en & mem_MPORT_455_mask) begin
      mem[mem_MPORT_455_addr] <= mem_MPORT_455_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_456_en & mem_MPORT_456_mask) begin
      mem[mem_MPORT_456_addr] <= mem_MPORT_456_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_457_en & mem_MPORT_457_mask) begin
      mem[mem_MPORT_457_addr] <= mem_MPORT_457_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_458_en & mem_MPORT_458_mask) begin
      mem[mem_MPORT_458_addr] <= mem_MPORT_458_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_459_en & mem_MPORT_459_mask) begin
      mem[mem_MPORT_459_addr] <= mem_MPORT_459_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_460_en & mem_MPORT_460_mask) begin
      mem[mem_MPORT_460_addr] <= mem_MPORT_460_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_461_en & mem_MPORT_461_mask) begin
      mem[mem_MPORT_461_addr] <= mem_MPORT_461_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_462_en & mem_MPORT_462_mask) begin
      mem[mem_MPORT_462_addr] <= mem_MPORT_462_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_463_en & mem_MPORT_463_mask) begin
      mem[mem_MPORT_463_addr] <= mem_MPORT_463_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_464_en & mem_MPORT_464_mask) begin
      mem[mem_MPORT_464_addr] <= mem_MPORT_464_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_465_en & mem_MPORT_465_mask) begin
      mem[mem_MPORT_465_addr] <= mem_MPORT_465_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_466_en & mem_MPORT_466_mask) begin
      mem[mem_MPORT_466_addr] <= mem_MPORT_466_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_467_en & mem_MPORT_467_mask) begin
      mem[mem_MPORT_467_addr] <= mem_MPORT_467_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_468_en & mem_MPORT_468_mask) begin
      mem[mem_MPORT_468_addr] <= mem_MPORT_468_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_469_en & mem_MPORT_469_mask) begin
      mem[mem_MPORT_469_addr] <= mem_MPORT_469_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_470_en & mem_MPORT_470_mask) begin
      mem[mem_MPORT_470_addr] <= mem_MPORT_470_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_471_en & mem_MPORT_471_mask) begin
      mem[mem_MPORT_471_addr] <= mem_MPORT_471_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_472_en & mem_MPORT_472_mask) begin
      mem[mem_MPORT_472_addr] <= mem_MPORT_472_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_473_en & mem_MPORT_473_mask) begin
      mem[mem_MPORT_473_addr] <= mem_MPORT_473_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_474_en & mem_MPORT_474_mask) begin
      mem[mem_MPORT_474_addr] <= mem_MPORT_474_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_475_en & mem_MPORT_475_mask) begin
      mem[mem_MPORT_475_addr] <= mem_MPORT_475_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_476_en & mem_MPORT_476_mask) begin
      mem[mem_MPORT_476_addr] <= mem_MPORT_476_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_477_en & mem_MPORT_477_mask) begin
      mem[mem_MPORT_477_addr] <= mem_MPORT_477_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_478_en & mem_MPORT_478_mask) begin
      mem[mem_MPORT_478_addr] <= mem_MPORT_478_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_479_en & mem_MPORT_479_mask) begin
      mem[mem_MPORT_479_addr] <= mem_MPORT_479_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_480_en & mem_MPORT_480_mask) begin
      mem[mem_MPORT_480_addr] <= mem_MPORT_480_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_481_en & mem_MPORT_481_mask) begin
      mem[mem_MPORT_481_addr] <= mem_MPORT_481_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_482_en & mem_MPORT_482_mask) begin
      mem[mem_MPORT_482_addr] <= mem_MPORT_482_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_483_en & mem_MPORT_483_mask) begin
      mem[mem_MPORT_483_addr] <= mem_MPORT_483_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_484_en & mem_MPORT_484_mask) begin
      mem[mem_MPORT_484_addr] <= mem_MPORT_484_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_485_en & mem_MPORT_485_mask) begin
      mem[mem_MPORT_485_addr] <= mem_MPORT_485_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_486_en & mem_MPORT_486_mask) begin
      mem[mem_MPORT_486_addr] <= mem_MPORT_486_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_487_en & mem_MPORT_487_mask) begin
      mem[mem_MPORT_487_addr] <= mem_MPORT_487_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_488_en & mem_MPORT_488_mask) begin
      mem[mem_MPORT_488_addr] <= mem_MPORT_488_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_489_en & mem_MPORT_489_mask) begin
      mem[mem_MPORT_489_addr] <= mem_MPORT_489_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_490_en & mem_MPORT_490_mask) begin
      mem[mem_MPORT_490_addr] <= mem_MPORT_490_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_491_en & mem_MPORT_491_mask) begin
      mem[mem_MPORT_491_addr] <= mem_MPORT_491_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_492_en & mem_MPORT_492_mask) begin
      mem[mem_MPORT_492_addr] <= mem_MPORT_492_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_493_en & mem_MPORT_493_mask) begin
      mem[mem_MPORT_493_addr] <= mem_MPORT_493_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_494_en & mem_MPORT_494_mask) begin
      mem[mem_MPORT_494_addr] <= mem_MPORT_494_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_495_en & mem_MPORT_495_mask) begin
      mem[mem_MPORT_495_addr] <= mem_MPORT_495_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_496_en & mem_MPORT_496_mask) begin
      mem[mem_MPORT_496_addr] <= mem_MPORT_496_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_497_en & mem_MPORT_497_mask) begin
      mem[mem_MPORT_497_addr] <= mem_MPORT_497_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_498_en & mem_MPORT_498_mask) begin
      mem[mem_MPORT_498_addr] <= mem_MPORT_498_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_499_en & mem_MPORT_499_mask) begin
      mem[mem_MPORT_499_addr] <= mem_MPORT_499_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_500_en & mem_MPORT_500_mask) begin
      mem[mem_MPORT_500_addr] <= mem_MPORT_500_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_501_en & mem_MPORT_501_mask) begin
      mem[mem_MPORT_501_addr] <= mem_MPORT_501_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_502_en & mem_MPORT_502_mask) begin
      mem[mem_MPORT_502_addr] <= mem_MPORT_502_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_503_en & mem_MPORT_503_mask) begin
      mem[mem_MPORT_503_addr] <= mem_MPORT_503_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_504_en & mem_MPORT_504_mask) begin
      mem[mem_MPORT_504_addr] <= mem_MPORT_504_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_505_en & mem_MPORT_505_mask) begin
      mem[mem_MPORT_505_addr] <= mem_MPORT_505_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_506_en & mem_MPORT_506_mask) begin
      mem[mem_MPORT_506_addr] <= mem_MPORT_506_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_507_en & mem_MPORT_507_mask) begin
      mem[mem_MPORT_507_addr] <= mem_MPORT_507_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_508_en & mem_MPORT_508_mask) begin
      mem[mem_MPORT_508_addr] <= mem_MPORT_508_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_509_en & mem_MPORT_509_mask) begin
      mem[mem_MPORT_509_addr] <= mem_MPORT_509_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_510_en & mem_MPORT_510_mask) begin
      mem[mem_MPORT_510_addr] <= mem_MPORT_510_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_511_en & mem_MPORT_511_mask) begin
      mem[mem_MPORT_511_addr] <= mem_MPORT_511_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_512_en & mem_MPORT_512_mask) begin
      mem[mem_MPORT_512_addr] <= mem_MPORT_512_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_15(
  input        clock,
  input        reset,
  input  [8:0] io_r_addr,
  output [1:0] io_r_data_0,
  output [1:0] io_r_data_1,
  output [1:0] io_r_data_2,
  output [1:0] io_r_data_3,
  input        io_w_en,
  input  [8:0] io_w_addr,
  input  [1:0] io_w_data_0,
  input  [1:0] io_w_data_1,
  input  [1:0] io_w_data_2,
  input  [1:0] io_w_data_3,
  input  [3:0] io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [8:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P_100 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P_100 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P_100 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P_100 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
endmodule
module MaxPeriodFibonacciLFSR_1(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  wire  _T_2 = state_7 ^ state_5 ^ state_4 ^ state_3; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T_2; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_4 <= state_3;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_5 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_5 <= state_4;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_6 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_6 <= state_5;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_7 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_7 <= state_6;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCacheDirectory_1(
  input         clock,
  input         reset,
  output        io_read_req_ready,
  input         io_read_req_valid,
  input  [31:0] io_read_req_bits_addr,
  output        io_read_resp_bits_hit,
  output [3:0]  io_read_resp_bits_chosenWay,
  output        io_read_resp_bits_isDirtyWay,
  output [18:0] io_read_resp_bits_tagRdVec_0,
  output [18:0] io_read_resp_bits_tagRdVec_1,
  output [18:0] io_read_resp_bits_tagRdVec_2,
  output [18:0] io_read_resp_bits_tagRdVec_3,
  output        io_write_req_ready,
  input         io_write_req_valid,
  input  [31:0] io_write_req_bits_addr,
  input  [3:0]  io_write_req_bits_way,
  input  [1:0]  io_write_req_bits_meta
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  tagArray_clock; // @[SRAM_1.scala 255:31]
  wire  tagArray_reset; // @[SRAM_1.scala 255:31]
  wire [8:0] tagArray_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [18:0] tagArray_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [18:0] tagArray_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [18:0] tagArray_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [18:0] tagArray_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  tagArray_io_w_en; // @[SRAM_1.scala 255:31]
  wire [8:0] tagArray_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [18:0] tagArray_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [18:0] tagArray_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [18:0] tagArray_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [18:0] tagArray_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] tagArray_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  metaArray_clock; // @[SRAM_1.scala 255:31]
  wire  metaArray_reset; // @[SRAM_1.scala 255:31]
  wire [8:0] metaArray_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  metaArray_io_w_en; // @[SRAM_1.scala 255:31]
  wire [8:0] metaArray_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] metaArray_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  replaceWay_lfsr_prng_clock; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_reset; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_7; // @[PRNG.scala 91:22]
  wire [8:0] rSet = io_read_req_bits_addr[12:4]; // @[Parameters.scala 50:11]
  wire [18:0] rTag = io_read_req_bits_addr[31:13]; // @[Parameters.scala 46:11]
  wire  ren = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  wire [8:0] wSet = io_write_req_bits_addr[12:4]; // @[Parameters.scala 50:11]
  wire [18:0] wTag = io_write_req_bits_addr[31:13]; // @[Parameters.scala 46:11]
  wire  wen = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _T_4 = io_write_req_bits_way[0] + io_write_req_bits_way[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_6 = io_write_req_bits_way[2] + io_write_req_bits_way[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_8 = _T_4 + _T_6; // @[Bitwise.scala 51:90]
  wire  _T_22 = ~reset; // @[Directory.scala 69:11]
  wire [18:0] rdata__0 = ren ? tagArray_io_r_data_0 : 19'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [18:0] rdata__1 = ren ? tagArray_io_r_data_1 : 19'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [18:0] rdata__2 = ren ? tagArray_io_r_data_2 : 19'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [18:0] rdata__3 = ren ? tagArray_io_r_data_3 : 19'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_0 = ren ? metaArray_io_r_data_0 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_1 = ren ? metaArray_io_r_data_1 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_2 = ren ? metaArray_io_r_data_2 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_3 = ren ? metaArray_io_r_data_3 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [7:0] _T_24 = {rdata_1_3,rdata_1_2,rdata_1_1,rdata_1_0}; // @[Directory.scala 82:52]
  wire  metaRdVec_0_valid = _T_24[0]; // @[Directory.scala 82:52]
  wire  metaRdVec_0_dirty = _T_24[1]; // @[Directory.scala 82:52]
  wire  metaRdVec_1_valid = _T_24[2]; // @[Directory.scala 82:52]
  wire  metaRdVec_1_dirty = _T_24[3]; // @[Directory.scala 82:52]
  wire  metaRdVec_2_valid = _T_24[4]; // @[Directory.scala 82:52]
  wire  metaRdVec_2_dirty = _T_24[5]; // @[Directory.scala 82:52]
  wire  metaRdVec_3_valid = _T_24[6]; // @[Directory.scala 82:52]
  wire  metaRdVec_3_dirty = _T_24[7]; // @[Directory.scala 82:52]
  wire  tagMatchVec_0 = rdata__0 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_1 = rdata__1 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_2 = rdata__2 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_3 = rdata__3 == rTag; // @[Directory.scala 85:46]
  wire  _matchWayOH_T = tagMatchVec_0 & metaRdVec_0_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_1 = tagMatchVec_1 & metaRdVec_1_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_2 = tagMatchVec_2 & metaRdVec_2_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_3 = tagMatchVec_3 & metaRdVec_3_valid; // @[Directory.scala 88:80]
  wire [3:0] matchWayOH = {_matchWayOH_T_3,_matchWayOH_T_2,_matchWayOH_T_1,_matchWayOH_T}; // @[Cat.scala 33:92]
  wire  invalidWayVec_0 = ~metaRdVec_0_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_1 = ~metaRdVec_1_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_2 = ~metaRdVec_2_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_3 = ~metaRdVec_3_valid; // @[Directory.scala 89:53]
  wire [3:0] _invalidWayOH_T_8 = invalidWayVec_2 ? 4'h4 : 4'h8; // @[Mux.scala 47:70]
  wire [3:0] _invalidWayOH_T_9 = invalidWayVec_1 ? 4'h2 : _invalidWayOH_T_8; // @[Mux.scala 47:70]
  wire [3:0] invalidWayOH = invalidWayVec_0 ? 4'h1 : _invalidWayOH_T_9; // @[Mux.scala 47:70]
  wire [3:0] _hasInvalidWay_T = {invalidWayVec_0,invalidWayVec_1,invalidWayVec_2,invalidWayVec_3}; // @[Cat.scala 33:92]
  wire  hasInvalidWay = |_hasInvalidWay_T; // @[Directory.scala 91:44]
  wire [7:0] replaceWay_lfsr = {replaceWay_lfsr_prng_io_out_7,replaceWay_lfsr_prng_io_out_6,
    replaceWay_lfsr_prng_io_out_5,replaceWay_lfsr_prng_io_out_4,replaceWay_lfsr_prng_io_out_3,
    replaceWay_lfsr_prng_io_out_2,replaceWay_lfsr_prng_io_out_1,replaceWay_lfsr_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [1:0] replaceWay_outputWay_shiftAmount = replaceWay_lfsr[1:0]; // @[DCache.scala 61:39]
  wire [3:0] replaceWay = 4'h1 << replaceWay_outputWay_shiftAmount; // @[OneHot.scala 64:12]
  wire  _replaceWayReg_T = ~io_read_req_valid; // @[Directory.scala 93:65]
  reg [3:0] replaceWayReg; // @[Reg.scala 19:16]
  wire  isHit = |matchWayOH; // @[Directory.scala 95:41]
  wire [3:0] _choseWayOH_T = hasInvalidWay ? invalidWayOH : replaceWayReg; // @[Directory.scala 96:51]
  wire [3:0] choseWayOH = isHit ? matchWayOH : _choseWayOH_T; // @[Directory.scala 96:28]
  wire [3:0] dirtyWayOH = {metaRdVec_3_dirty,metaRdVec_2_dirty,metaRdVec_1_dirty,metaRdVec_0_dirty}; // @[Cat.scala 33:92]
  wire [3:0] _isDirtyWay_T = choseWayOH & dirtyWayOH; // @[Directory.scala 98:38]
  wire [1:0] _T_37 = choseWayOH[0] + choseWayOH[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_39 = choseWayOH[2] + choseWayOH[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_41 = _T_37 + _T_39; // @[Bitwise.scala 51:90]
  SRAMArray_2P_14 tagArray ( // @[SRAM_1.scala 255:31]
    .clock(tagArray_clock),
    .reset(tagArray_reset),
    .io_r_addr(tagArray_io_r_addr),
    .io_r_data_0(tagArray_io_r_data_0),
    .io_r_data_1(tagArray_io_r_data_1),
    .io_r_data_2(tagArray_io_r_data_2),
    .io_r_data_3(tagArray_io_r_data_3),
    .io_w_en(tagArray_io_w_en),
    .io_w_addr(tagArray_io_w_addr),
    .io_w_data_0(tagArray_io_w_data_0),
    .io_w_data_1(tagArray_io_w_data_1),
    .io_w_data_2(tagArray_io_w_data_2),
    .io_w_data_3(tagArray_io_w_data_3),
    .io_w_maskOH(tagArray_io_w_maskOH)
  );
  SRAMArray_2P_15 metaArray ( // @[SRAM_1.scala 255:31]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_addr(metaArray_io_r_addr),
    .io_r_data_0(metaArray_io_r_data_0),
    .io_r_data_1(metaArray_io_r_data_1),
    .io_r_data_2(metaArray_io_r_data_2),
    .io_r_data_3(metaArray_io_r_data_3),
    .io_w_en(metaArray_io_w_en),
    .io_w_addr(metaArray_io_w_addr),
    .io_w_data_0(metaArray_io_w_data_0),
    .io_w_data_1(metaArray_io_w_data_1),
    .io_w_data_2(metaArray_io_w_data_2),
    .io_w_data_3(metaArray_io_w_data_3),
    .io_w_maskOH(metaArray_io_w_maskOH)
  );
  MaxPeriodFibonacciLFSR_1 replaceWay_lfsr_prng ( // @[PRNG.scala 91:22]
    .clock(replaceWay_lfsr_prng_clock),
    .reset(replaceWay_lfsr_prng_reset),
    .io_out_0(replaceWay_lfsr_prng_io_out_0),
    .io_out_1(replaceWay_lfsr_prng_io_out_1),
    .io_out_2(replaceWay_lfsr_prng_io_out_2),
    .io_out_3(replaceWay_lfsr_prng_io_out_3),
    .io_out_4(replaceWay_lfsr_prng_io_out_4),
    .io_out_5(replaceWay_lfsr_prng_io_out_5),
    .io_out_6(replaceWay_lfsr_prng_io_out_6),
    .io_out_7(replaceWay_lfsr_prng_io_out_7)
  );
  assign io_read_req_ready = 1'h1; // @[Directory.scala 75:29]
  assign io_read_resp_bits_hit = |matchWayOH; // @[Directory.scala 95:41]
  assign io_read_resp_bits_chosenWay = isHit ? matchWayOH : _choseWayOH_T; // @[Directory.scala 96:28]
  assign io_read_resp_bits_isDirtyWay = |_isDirtyWay_T; // @[Directory.scala 98:53]
  assign io_read_resp_bits_tagRdVec_0 = ren ? tagArray_io_r_data_0 : 19'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_1 = ren ? tagArray_io_r_data_1 : 19'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_2 = ren ? tagArray_io_r_data_2 : 19'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_3 = ren ? tagArray_io_r_data_3 : 19'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_write_req_ready = 1'h1; // @[Directory.scala 76:29]
  assign tagArray_clock = clock;
  assign tagArray_reset = reset;
  assign tagArray_io_r_addr = rSet; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign tagArray_io_w_en = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  assign tagArray_io_w_addr = wSet; // @[Directory.scala 112:15 SRAM_1.scala 237:19]
  assign tagArray_io_w_data_0 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_1 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_2 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_3 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_maskOH = io_write_req_bits_way; // @[Directory.scala 112:15 SRAM_1.scala 239:21]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r_addr = rSet; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign metaArray_io_w_en = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  assign metaArray_io_w_addr = wSet; // @[Directory.scala 112:15 SRAM_1.scala 237:19]
  assign metaArray_io_w_data_0 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_1 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_2 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_3 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_maskOH = io_write_req_bits_way; // @[Directory.scala 112:15 SRAM_1.scala 239:21]
  assign replaceWay_lfsr_prng_clock = clock;
  assign replaceWay_lfsr_prng_reset = reset;
  always @(posedge clock) begin
    if (_replaceWayReg_T) begin // @[Reg.scala 20:18]
      replaceWayReg <= replaceWay; // @[Reg.scala 20:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_8 < 3'h2)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Error directory write way has multiple valid bit! ==>%d\n    at Directory.scala:69 assert(PopCount(wWay) < 2.U, cf\"Error directory write way has multiple valid bit! ==>${PopCount(wWay)}\")\n"
            ,_T_8); // @[Directory.scala 69:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_8 < 3'h2) & ~reset) begin
          $fatal; // @[Directory.scala 69:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & ~(_T_41 == 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Error chosenWay has multiple valid bit!\n    at Directory.scala:101 assert(PopCount(choseWayOH) === 1.U, \"Error chosenWay has multiple valid bit!\")\n"
            ); // @[Directory.scala 101:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_41 == 3'h1) & _T_22) begin
          $fatal; // @[Directory.scala 101:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wen & _T_22 & ~(_T_8 <= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: write error, tring to write multiple ways\n    at SRAM_1.scala:235 assert(PopCount(mask) <= 1.U, \"write error, tring to write multiple ways\")\n"
            ); // @[SRAM_1.scala 235:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_8 <= 3'h1) & (wen & _T_22)) begin
          $fatal; // @[SRAM_1.scala 235:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wen & _T_22 & ~(_T_8 <= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: write error, tring to write multiple ways\n    at SRAM_1.scala:235 assert(PopCount(mask) <= 1.U, \"write error, tring to write multiple ways\")\n"
            ); // @[SRAM_1.scala 235:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_8 <= 3'h1) & (wen & _T_22)) begin
          $fatal; // @[SRAM_1.scala 235:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  replaceWayReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_1(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input         io_in_0_bits_dirInfo_hit,
  input  [3:0]  io_in_0_bits_dirInfo_chosenWay,
  input         io_in_0_bits_dirInfo_isDirtyWay,
  input  [18:0] io_in_0_bits_dirtyTag,
  input  [31:0] io_in_0_bits_data_0,
  input  [31:0] io_in_0_bits_data_1,
  input  [31:0] io_in_0_bits_data_2,
  input  [31:0] io_in_0_bits_data_3,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input         io_in_1_bits_dirInfo_hit,
  input  [3:0]  io_in_1_bits_dirInfo_chosenWay,
  input         io_in_1_bits_dirInfo_isDirtyWay,
  input  [18:0] io_in_1_bits_dirtyTag,
  input  [31:0] io_in_1_bits_data_0,
  input  [31:0] io_in_1_bits_data_1,
  input  [31:0] io_in_1_bits_data_2,
  input  [31:0] io_in_1_bits_data_3,
  input  [31:0] io_in_1_bits_storeData,
  input  [3:0]  io_in_1_bits_storeMask,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output        io_out_bits_dirInfo_hit,
  output [3:0]  io_out_bits_dirInfo_chosenWay,
  output        io_out_bits_dirInfo_isDirtyWay,
  output [18:0] io_out_bits_dirtyTag,
  output [31:0] io_out_bits_data_0,
  output [31:0] io_out_bits_data_1,
  output [31:0] io_out_bits_data_2,
  output [31:0] io_out_bits_data_3,
  output        io_out_bits_isStore,
  output [31:0] io_out_bits_storeData,
  output [3:0]  io_out_bits_storeMask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_dirInfo_hit = io_in_0_valid ? io_in_0_bits_dirInfo_hit : io_in_1_bits_dirInfo_hit; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_dirInfo_chosenWay = io_in_0_valid ? io_in_0_bits_dirInfo_chosenWay : io_in_1_bits_dirInfo_chosenWay
    ; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_dirInfo_isDirtyWay = io_in_0_valid ? io_in_0_bits_dirInfo_isDirtyWay :
    io_in_1_bits_dirInfo_isDirtyWay; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_dirtyTag = io_in_0_valid ? io_in_0_bits_dirtyTag : io_in_1_bits_dirtyTag; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data_0 = io_in_0_valid ? io_in_0_bits_data_0 : io_in_1_bits_data_0; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data_1 = io_in_0_valid ? io_in_0_bits_data_1 : io_in_1_bits_data_1; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data_2 = io_in_0_valid ? io_in_0_bits_data_2 : io_in_1_bits_data_2; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data_3 = io_in_0_valid ? io_in_0_bits_data_3 : io_in_1_bits_data_3; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_isStore = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_storeData = io_in_0_valid ? 32'h0 : io_in_1_bits_storeData; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_storeMask = io_in_0_valid ? 4'h0 : io_in_1_bits_storeMask; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_2(
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [31:0]  io_in_0_bits_address,
  input  [127:0] io_in_0_bits_data,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [31:0]  io_in_1_bits_address,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_opcode,
  output [31:0]  io_out_bits_address,
  output [127:0] io_out_bits_data
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_opcode = io_in_0_valid ? 3'h2 : 3'h4; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_address = io_in_0_valid ? io_in_0_bits_address : io_in_1_bits_address; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : 128'h0; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_3(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_data,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_data
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_4(
  output  io_in_0_ready,
  input   io_in_0_valid,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input   io_out_ready,
  output  io_out_valid
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
endmodule
module Arbiter_5(
  input        io_in_0_valid,
  input  [8:0] io_in_0_bits_set,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [8:0] io_in_1_bits_set,
  output       io_out_valid,
  output [8:0] io_out_bits_set
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_set = io_in_0_valid ? io_in_0_bits_set : io_in_1_bits_set; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_6(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  output        io_out_valid,
  output [31:0] io_out_bits_addr
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_7(
  input         io_in_0_valid,
  input  [8:0]  io_in_0_bits_set,
  input  [31:0] io_in_0_bits_data_0,
  input  [31:0] io_in_0_bits_data_1,
  input  [31:0] io_in_0_bits_data_2,
  input  [31:0] io_in_0_bits_data_3,
  input  [3:0]  io_in_0_bits_blockMask,
  input  [3:0]  io_in_0_bits_way,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [8:0]  io_in_1_bits_set,
  input  [31:0] io_in_1_bits_data_0,
  input  [31:0] io_in_1_bits_data_1,
  input  [31:0] io_in_1_bits_data_2,
  input  [31:0] io_in_1_bits_data_3,
  input  [3:0]  io_in_1_bits_way,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [8:0]  io_in_2_bits_set,
  input  [31:0] io_in_2_bits_data_0,
  input  [31:0] io_in_2_bits_data_1,
  input  [31:0] io_in_2_bits_data_2,
  input  [31:0] io_in_2_bits_data_3,
  input  [3:0]  io_in_2_bits_blockMask,
  input  [3:0]  io_in_2_bits_way,
  output        io_out_valid,
  output [8:0]  io_out_bits_set,
  output [31:0] io_out_bits_data_0,
  output [31:0] io_out_bits_data_1,
  output [31:0] io_out_bits_data_2,
  output [31:0] io_out_bits_data_3,
  output [3:0]  io_out_bits_blockMask,
  output [3:0]  io_out_bits_way
);
  wire [8:0] _GEN_1 = io_in_1_valid ? io_in_1_bits_set : io_in_2_bits_set; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [31:0] _GEN_3 = io_in_1_valid ? io_in_1_bits_data_0 : io_in_2_bits_data_0; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [31:0] _GEN_4 = io_in_1_valid ? io_in_1_bits_data_1 : io_in_2_bits_data_1; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [31:0] _GEN_5 = io_in_1_valid ? io_in_1_bits_data_2 : io_in_2_bits_data_2; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [31:0] _GEN_6 = io_in_1_valid ? io_in_1_bits_data_3 : io_in_2_bits_data_3; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [3:0] _GEN_7 = io_in_1_valid ? 4'hf : io_in_2_bits_blockMask; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [3:0] _GEN_8 = io_in_1_valid ? io_in_1_bits_way : io_in_2_bits_way; // @[Arbiter.scala 136:15 138:26 140:19]
  wire  grant_2 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_2_ready = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_2 | io_in_2_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_set = io_in_0_valid ? io_in_0_bits_set : _GEN_1; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_data_0 = io_in_0_valid ? io_in_0_bits_data_0 : _GEN_3; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_data_1 = io_in_0_valid ? io_in_0_bits_data_1 : _GEN_4; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_data_2 = io_in_0_valid ? io_in_0_bits_data_2 : _GEN_5; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_data_3 = io_in_0_valid ? io_in_0_bits_data_3 : _GEN_6; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_blockMask = io_in_0_valid ? io_in_0_bits_blockMask : _GEN_7; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_way = io_in_0_valid ? io_in_0_bits_way : _GEN_8; // @[Arbiter.scala 138:26 140:19]
endmodule
module Arbiter_8(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [3:0]  io_in_0_bits_way,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [3:0]  io_in_1_bits_way,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input  [3:0]  io_in_2_bits_way,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [3:0]  io_out_bits_way,
  output [1:0]  io_out_bits_meta
);
  wire [31:0] _GEN_1 = io_in_1_valid ? io_in_1_bits_addr : io_in_2_bits_addr; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [3:0] _GEN_2 = io_in_1_valid ? io_in_1_bits_way : io_in_2_bits_way; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [1:0] _GEN_3 = io_in_1_valid ? 2'h1 : 2'h3; // @[Arbiter.scala 136:15 138:26 140:19]
  wire  grant_2 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_2_ready = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_2 | io_in_2_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_1; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_way = io_in_0_valid ? io_in_0_bits_way : _GEN_2; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_meta = io_in_0_valid ? 2'h3 : _GEN_3; // @[Arbiter.scala 138:26 140:19]
endmodule
module DCache(
  input          clock,
  input          reset,
  output         io_read_req_ready,
  input          io_read_req_valid,
  input  [31:0]  io_read_req_bits_addr,
  input          io_read_resp_ready,
  output         io_read_resp_valid,
  output [31:0]  io_read_resp_bits_data,
  output         io_write_req_ready,
  input          io_write_req_valid,
  input  [31:0]  io_write_req_bits_addr,
  input  [31:0]  io_write_req_bits_data,
  input  [3:0]   io_write_req_bits_mask,
  input          io_write_resp_ready,
  output         io_write_resp_valid,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [2:0]   io_tlbus_req_bits_opcode,
  output [31:0]  io_tlbus_req_bits_address,
  output [127:0] io_tlbus_req_bits_data,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data,
  input          io_flush
);
  wire  loadPipe_clock; // @[DCache.scala 82:26]
  wire  loadPipe_reset; // @[DCache.scala 82:26]
  wire  loadPipe_io_load_req_ready; // @[DCache.scala 82:26]
  wire  loadPipe_io_load_req_valid; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_load_req_bits_addr; // @[DCache.scala 82:26]
  wire  loadPipe_io_load_resp_ready; // @[DCache.scala 82:26]
  wire  loadPipe_io_load_resp_valid; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_load_resp_bits_data; // @[DCache.scala 82:26]
  wire  loadPipe_io_dir_req_ready; // @[DCache.scala 82:26]
  wire  loadPipe_io_dir_req_valid; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dir_req_bits_addr; // @[DCache.scala 82:26]
  wire  loadPipe_io_dir_resp_bits_hit; // @[DCache.scala 82:26]
  wire [3:0] loadPipe_io_dir_resp_bits_chosenWay; // @[DCache.scala 82:26]
  wire  loadPipe_io_dir_resp_bits_isDirtyWay; // @[DCache.scala 82:26]
  wire [18:0] loadPipe_io_dir_resp_bits_tagRdVec_0; // @[DCache.scala 82:26]
  wire [18:0] loadPipe_io_dir_resp_bits_tagRdVec_1; // @[DCache.scala 82:26]
  wire [18:0] loadPipe_io_dir_resp_bits_tagRdVec_2; // @[DCache.scala 82:26]
  wire [18:0] loadPipe_io_dir_resp_bits_tagRdVec_3; // @[DCache.scala 82:26]
  wire  loadPipe_io_dataBank_req_ready; // @[DCache.scala 82:26]
  wire  loadPipe_io_dataBank_req_valid; // @[DCache.scala 82:26]
  wire [8:0] loadPipe_io_dataBank_req_bits_set; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_0_0; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_0_1; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_0_2; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_0_3; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_1_0; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_1_1; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_1_2; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_1_3; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_2_0; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_2_1; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_2_2; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_2_3; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_3_0; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_3_1; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_3_2; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_dataBank_resp_3_3; // @[DCache.scala 82:26]
  wire  loadPipe_io_mshr_ready; // @[DCache.scala 82:26]
  wire  loadPipe_io_mshr_valid; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_mshr_bits_addr; // @[DCache.scala 82:26]
  wire  loadPipe_io_mshr_bits_dirInfo_hit; // @[DCache.scala 82:26]
  wire [3:0] loadPipe_io_mshr_bits_dirInfo_chosenWay; // @[DCache.scala 82:26]
  wire  loadPipe_io_mshr_bits_dirInfo_isDirtyWay; // @[DCache.scala 82:26]
  wire [18:0] loadPipe_io_mshr_bits_dirtyTag; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_mshr_bits_data_0; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_mshr_bits_data_1; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_mshr_bits_data_2; // @[DCache.scala 82:26]
  wire [31:0] loadPipe_io_mshr_bits_data_3; // @[DCache.scala 82:26]
  wire  storePipe_clock; // @[DCache.scala 83:27]
  wire  storePipe_reset; // @[DCache.scala 83:27]
  wire  storePipe_io_store_req_ready; // @[DCache.scala 83:27]
  wire  storePipe_io_store_req_valid; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_store_req_bits_addr; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_store_req_bits_data; // @[DCache.scala 83:27]
  wire [3:0] storePipe_io_store_req_bits_mask; // @[DCache.scala 83:27]
  wire  storePipe_io_store_resp_ready; // @[DCache.scala 83:27]
  wire  storePipe_io_store_resp_valid; // @[DCache.scala 83:27]
  wire  storePipe_io_dir_read_req_valid; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dir_read_req_bits_addr; // @[DCache.scala 83:27]
  wire  storePipe_io_dir_read_resp_bits_hit; // @[DCache.scala 83:27]
  wire [3:0] storePipe_io_dir_read_resp_bits_chosenWay; // @[DCache.scala 83:27]
  wire  storePipe_io_dir_read_resp_bits_isDirtyWay; // @[DCache.scala 83:27]
  wire [18:0] storePipe_io_dir_read_resp_bits_tagRdVec_0; // @[DCache.scala 83:27]
  wire [18:0] storePipe_io_dir_read_resp_bits_tagRdVec_1; // @[DCache.scala 83:27]
  wire [18:0] storePipe_io_dir_read_resp_bits_tagRdVec_2; // @[DCache.scala 83:27]
  wire [18:0] storePipe_io_dir_read_resp_bits_tagRdVec_3; // @[DCache.scala 83:27]
  wire  storePipe_io_dir_write_req_valid; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dir_write_req_bits_addr; // @[DCache.scala 83:27]
  wire [3:0] storePipe_io_dir_write_req_bits_way; // @[DCache.scala 83:27]
  wire  storePipe_io_dataBank_read_req_valid; // @[DCache.scala 83:27]
  wire [8:0] storePipe_io_dataBank_read_req_bits_set; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_0_0; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_0_1; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_0_2; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_0_3; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_1_0; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_1_1; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_1_2; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_1_3; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_2_0; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_2_1; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_2_2; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_2_3; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_3_0; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_3_1; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_3_2; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_read_resp_3_3; // @[DCache.scala 83:27]
  wire  storePipe_io_dataBank_write_req_valid; // @[DCache.scala 83:27]
  wire [8:0] storePipe_io_dataBank_write_req_bits_set; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_write_req_bits_data_0; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_write_req_bits_data_1; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_write_req_bits_data_2; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_dataBank_write_req_bits_data_3; // @[DCache.scala 83:27]
  wire [3:0] storePipe_io_dataBank_write_req_bits_blockMask; // @[DCache.scala 83:27]
  wire [3:0] storePipe_io_dataBank_write_req_bits_way; // @[DCache.scala 83:27]
  wire  storePipe_io_mshr_ready; // @[DCache.scala 83:27]
  wire  storePipe_io_mshr_valid; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_mshr_bits_addr; // @[DCache.scala 83:27]
  wire  storePipe_io_mshr_bits_dirInfo_hit; // @[DCache.scala 83:27]
  wire [3:0] storePipe_io_mshr_bits_dirInfo_chosenWay; // @[DCache.scala 83:27]
  wire  storePipe_io_mshr_bits_dirInfo_isDirtyWay; // @[DCache.scala 83:27]
  wire [18:0] storePipe_io_mshr_bits_dirtyTag; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_mshr_bits_data_0; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_mshr_bits_data_1; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_mshr_bits_data_2; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_mshr_bits_data_3; // @[DCache.scala 83:27]
  wire [31:0] storePipe_io_mshr_bits_storeData; // @[DCache.scala 83:27]
  wire [3:0] storePipe_io_mshr_bits_storeMask; // @[DCache.scala 83:27]
  wire  storePipe_io_flush; // @[DCache.scala 83:27]
  wire  mshr_clock; // @[DCache.scala 84:22]
  wire  mshr_reset; // @[DCache.scala 84:22]
  wire  mshr_io_req_ready; // @[DCache.scala 84:22]
  wire  mshr_io_req_valid; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_req_bits_addr; // @[DCache.scala 84:22]
  wire  mshr_io_req_bits_dirInfo_hit; // @[DCache.scala 84:22]
  wire [3:0] mshr_io_req_bits_dirInfo_chosenWay; // @[DCache.scala 84:22]
  wire  mshr_io_req_bits_dirInfo_isDirtyWay; // @[DCache.scala 84:22]
  wire [18:0] mshr_io_req_bits_dirtyTag; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_req_bits_data_0; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_req_bits_data_1; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_req_bits_data_2; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_req_bits_data_3; // @[DCache.scala 84:22]
  wire  mshr_io_req_bits_isStore; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_req_bits_storeData; // @[DCache.scala 84:22]
  wire [3:0] mshr_io_req_bits_storeMask; // @[DCache.scala 84:22]
  wire  mshr_io_resp_load_ready; // @[DCache.scala 84:22]
  wire  mshr_io_resp_load_valid; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_resp_load_bits_data; // @[DCache.scala 84:22]
  wire  mshr_io_resp_store_ready; // @[DCache.scala 84:22]
  wire  mshr_io_resp_store_valid; // @[DCache.scala 84:22]
  wire  mshr_io_tasks_refill_req_valid; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_tasks_refill_req_bits_addr; // @[DCache.scala 84:22]
  wire [3:0] mshr_io_tasks_refill_req_bits_chosenWay; // @[DCache.scala 84:22]
  wire  mshr_io_tasks_refill_resp_ready; // @[DCache.scala 84:22]
  wire  mshr_io_tasks_refill_resp_valid; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_tasks_refill_resp_bits_data; // @[DCache.scala 84:22]
  wire  mshr_io_tasks_writeback_req_valid; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_addr; // @[DCache.scala 84:22]
  wire [18:0] mshr_io_tasks_writeback_req_bits_dirtyTag; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_data_0; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_data_1; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_data_2; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_data_3; // @[DCache.scala 84:22]
  wire  mshr_io_tasks_writeback_resp_ready; // @[DCache.scala 84:22]
  wire  mshr_io_tasks_writeback_resp_valid; // @[DCache.scala 84:22]
  wire  mshr_io_dirWrite_req_ready; // @[DCache.scala 84:22]
  wire  mshr_io_dirWrite_req_valid; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_dirWrite_req_bits_addr; // @[DCache.scala 84:22]
  wire [3:0] mshr_io_dirWrite_req_bits_way; // @[DCache.scala 84:22]
  wire  mshr_io_dataWrite_req_ready; // @[DCache.scala 84:22]
  wire  mshr_io_dataWrite_req_valid; // @[DCache.scala 84:22]
  wire [8:0] mshr_io_dataWrite_req_bits_set; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_dataWrite_req_bits_data_0; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_dataWrite_req_bits_data_1; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_dataWrite_req_bits_data_2; // @[DCache.scala 84:22]
  wire [31:0] mshr_io_dataWrite_req_bits_data_3; // @[DCache.scala 84:22]
  wire [3:0] mshr_io_dataWrite_req_bits_blockMask; // @[DCache.scala 84:22]
  wire [3:0] mshr_io_dataWrite_req_bits_way; // @[DCache.scala 84:22]
  wire  mshr_io_flush; // @[DCache.scala 84:22]
  wire  refillPipe_clock; // @[DCache.scala 85:28]
  wire  refillPipe_reset; // @[DCache.scala 85:28]
  wire  refillPipe_io_req_ready; // @[DCache.scala 85:28]
  wire  refillPipe_io_req_valid; // @[DCache.scala 85:28]
  wire [31:0] refillPipe_io_req_bits_addr; // @[DCache.scala 85:28]
  wire [3:0] refillPipe_io_req_bits_chosenWay; // @[DCache.scala 85:28]
  wire  refillPipe_io_resp_valid; // @[DCache.scala 85:28]
  wire [31:0] refillPipe_io_resp_bits_data; // @[DCache.scala 85:28]
  wire  refillPipe_io_tlbus_req_ready; // @[DCache.scala 85:28]
  wire  refillPipe_io_tlbus_req_valid; // @[DCache.scala 85:28]
  wire [31:0] refillPipe_io_tlbus_req_bits_address; // @[DCache.scala 85:28]
  wire  refillPipe_io_tlbus_resp_ready; // @[DCache.scala 85:28]
  wire  refillPipe_io_tlbus_resp_valid; // @[DCache.scala 85:28]
  wire [2:0] refillPipe_io_tlbus_resp_bits_opcode; // @[DCache.scala 85:28]
  wire [127:0] refillPipe_io_tlbus_resp_bits_data; // @[DCache.scala 85:28]
  wire  refillPipe_io_dirWrite_req_ready; // @[DCache.scala 85:28]
  wire  refillPipe_io_dirWrite_req_valid; // @[DCache.scala 85:28]
  wire [31:0] refillPipe_io_dirWrite_req_bits_addr; // @[DCache.scala 85:28]
  wire [3:0] refillPipe_io_dirWrite_req_bits_way; // @[DCache.scala 85:28]
  wire  refillPipe_io_dataWrite_req_ready; // @[DCache.scala 85:28]
  wire  refillPipe_io_dataWrite_req_valid; // @[DCache.scala 85:28]
  wire [8:0] refillPipe_io_dataWrite_req_bits_set; // @[DCache.scala 85:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_0; // @[DCache.scala 85:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_1; // @[DCache.scala 85:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_2; // @[DCache.scala 85:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_3; // @[DCache.scala 85:28]
  wire [3:0] refillPipe_io_dataWrite_req_bits_way; // @[DCache.scala 85:28]
  wire  wb_clock; // @[DCache.scala 86:20]
  wire  wb_reset; // @[DCache.scala 86:20]
  wire  wb_io_req_ready; // @[DCache.scala 86:20]
  wire  wb_io_req_valid; // @[DCache.scala 86:20]
  wire [31:0] wb_io_req_bits_addr; // @[DCache.scala 86:20]
  wire [18:0] wb_io_req_bits_dirtyTag; // @[DCache.scala 86:20]
  wire [31:0] wb_io_req_bits_data_0; // @[DCache.scala 86:20]
  wire [31:0] wb_io_req_bits_data_1; // @[DCache.scala 86:20]
  wire [31:0] wb_io_req_bits_data_2; // @[DCache.scala 86:20]
  wire [31:0] wb_io_req_bits_data_3; // @[DCache.scala 86:20]
  wire  wb_io_resp_valid; // @[DCache.scala 86:20]
  wire  wb_io_tlbus_req_ready; // @[DCache.scala 86:20]
  wire  wb_io_tlbus_req_valid; // @[DCache.scala 86:20]
  wire [31:0] wb_io_tlbus_req_bits_address; // @[DCache.scala 86:20]
  wire [127:0] wb_io_tlbus_req_bits_data; // @[DCache.scala 86:20]
  wire  wb_io_tlbus_resp_ready; // @[DCache.scala 86:20]
  wire  wb_io_tlbus_resp_valid; // @[DCache.scala 86:20]
  wire  db_clock; // @[DCache.scala 87:20]
  wire  db_reset; // @[DCache.scala 87:20]
  wire  db_io_read_req_ready; // @[DCache.scala 87:20]
  wire  db_io_read_req_valid; // @[DCache.scala 87:20]
  wire [8:0] db_io_read_req_bits_set; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_0_0; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_0_1; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_0_2; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_0_3; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_1_0; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_1_1; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_1_2; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_1_3; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_2_0; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_2_1; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_2_2; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_2_3; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_3_0; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_3_1; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_3_2; // @[DCache.scala 87:20]
  wire [31:0] db_io_read_resp_3_3; // @[DCache.scala 87:20]
  wire  db_io_write_req_ready; // @[DCache.scala 87:20]
  wire  db_io_write_req_valid; // @[DCache.scala 87:20]
  wire [8:0] db_io_write_req_bits_set; // @[DCache.scala 87:20]
  wire [31:0] db_io_write_req_bits_data_0; // @[DCache.scala 87:20]
  wire [31:0] db_io_write_req_bits_data_1; // @[DCache.scala 87:20]
  wire [31:0] db_io_write_req_bits_data_2; // @[DCache.scala 87:20]
  wire [31:0] db_io_write_req_bits_data_3; // @[DCache.scala 87:20]
  wire [3:0] db_io_write_req_bits_blockMask; // @[DCache.scala 87:20]
  wire [3:0] db_io_write_req_bits_way; // @[DCache.scala 87:20]
  wire  dir_clock; // @[DCache.scala 88:21]
  wire  dir_reset; // @[DCache.scala 88:21]
  wire  dir_io_read_req_ready; // @[DCache.scala 88:21]
  wire  dir_io_read_req_valid; // @[DCache.scala 88:21]
  wire [31:0] dir_io_read_req_bits_addr; // @[DCache.scala 88:21]
  wire  dir_io_read_resp_bits_hit; // @[DCache.scala 88:21]
  wire [3:0] dir_io_read_resp_bits_chosenWay; // @[DCache.scala 88:21]
  wire  dir_io_read_resp_bits_isDirtyWay; // @[DCache.scala 88:21]
  wire [18:0] dir_io_read_resp_bits_tagRdVec_0; // @[DCache.scala 88:21]
  wire [18:0] dir_io_read_resp_bits_tagRdVec_1; // @[DCache.scala 88:21]
  wire [18:0] dir_io_read_resp_bits_tagRdVec_2; // @[DCache.scala 88:21]
  wire [18:0] dir_io_read_resp_bits_tagRdVec_3; // @[DCache.scala 88:21]
  wire  dir_io_write_req_ready; // @[DCache.scala 88:21]
  wire  dir_io_write_req_valid; // @[DCache.scala 88:21]
  wire [31:0] dir_io_write_req_bits_addr; // @[DCache.scala 88:21]
  wire [3:0] dir_io_write_req_bits_way; // @[DCache.scala 88:21]
  wire [1:0] dir_io_write_req_bits_meta; // @[DCache.scala 88:21]
  wire  mshrReqArb_io_in_0_ready; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_in_0_valid; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_0_bits_addr; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_in_0_bits_dirInfo_hit; // @[DCache.scala 109:28]
  wire [3:0] mshrReqArb_io_in_0_bits_dirInfo_chosenWay; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_in_0_bits_dirInfo_isDirtyWay; // @[DCache.scala 109:28]
  wire [18:0] mshrReqArb_io_in_0_bits_dirtyTag; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_0_bits_data_0; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_0_bits_data_1; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_0_bits_data_2; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_0_bits_data_3; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_in_1_ready; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_in_1_valid; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_1_bits_addr; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_in_1_bits_dirInfo_hit; // @[DCache.scala 109:28]
  wire [3:0] mshrReqArb_io_in_1_bits_dirInfo_chosenWay; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_in_1_bits_dirInfo_isDirtyWay; // @[DCache.scala 109:28]
  wire [18:0] mshrReqArb_io_in_1_bits_dirtyTag; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_1_bits_data_0; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_1_bits_data_1; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_1_bits_data_2; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_1_bits_data_3; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_in_1_bits_storeData; // @[DCache.scala 109:28]
  wire [3:0] mshrReqArb_io_in_1_bits_storeMask; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_out_ready; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_out_valid; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_out_bits_addr; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_out_bits_dirInfo_hit; // @[DCache.scala 109:28]
  wire [3:0] mshrReqArb_io_out_bits_dirInfo_chosenWay; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_out_bits_dirInfo_isDirtyWay; // @[DCache.scala 109:28]
  wire [18:0] mshrReqArb_io_out_bits_dirtyTag; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_out_bits_data_0; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_out_bits_data_1; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_out_bits_data_2; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_out_bits_data_3; // @[DCache.scala 109:28]
  wire  mshrReqArb_io_out_bits_isStore; // @[DCache.scala 109:28]
  wire [31:0] mshrReqArb_io_out_bits_storeData; // @[DCache.scala 109:28]
  wire [3:0] mshrReqArb_io_out_bits_storeMask; // @[DCache.scala 109:28]
  wire  tlbusReqArb_io_in_0_ready; // @[DCache.scala 114:29]
  wire  tlbusReqArb_io_in_0_valid; // @[DCache.scala 114:29]
  wire [31:0] tlbusReqArb_io_in_0_bits_address; // @[DCache.scala 114:29]
  wire [127:0] tlbusReqArb_io_in_0_bits_data; // @[DCache.scala 114:29]
  wire  tlbusReqArb_io_in_1_ready; // @[DCache.scala 114:29]
  wire  tlbusReqArb_io_in_1_valid; // @[DCache.scala 114:29]
  wire [31:0] tlbusReqArb_io_in_1_bits_address; // @[DCache.scala 114:29]
  wire  tlbusReqArb_io_out_ready; // @[DCache.scala 114:29]
  wire  tlbusReqArb_io_out_valid; // @[DCache.scala 114:29]
  wire [2:0] tlbusReqArb_io_out_bits_opcode; // @[DCache.scala 114:29]
  wire [31:0] tlbusReqArb_io_out_bits_address; // @[DCache.scala 114:29]
  wire [127:0] tlbusReqArb_io_out_bits_data; // @[DCache.scala 114:29]
  wire  loadRespArb_io_in_0_ready; // @[DCache.scala 126:29]
  wire  loadRespArb_io_in_0_valid; // @[DCache.scala 126:29]
  wire [31:0] loadRespArb_io_in_0_bits_data; // @[DCache.scala 126:29]
  wire  loadRespArb_io_in_1_ready; // @[DCache.scala 126:29]
  wire  loadRespArb_io_in_1_valid; // @[DCache.scala 126:29]
  wire [31:0] loadRespArb_io_in_1_bits_data; // @[DCache.scala 126:29]
  wire  loadRespArb_io_out_ready; // @[DCache.scala 126:29]
  wire  loadRespArb_io_out_valid; // @[DCache.scala 126:29]
  wire [31:0] loadRespArb_io_out_bits_data; // @[DCache.scala 126:29]
  wire  storeRespArb_io_in_0_ready; // @[DCache.scala 131:30]
  wire  storeRespArb_io_in_0_valid; // @[DCache.scala 131:30]
  wire  storeRespArb_io_in_1_ready; // @[DCache.scala 131:30]
  wire  storeRespArb_io_in_1_valid; // @[DCache.scala 131:30]
  wire  storeRespArb_io_out_ready; // @[DCache.scala 131:30]
  wire  storeRespArb_io_out_valid; // @[DCache.scala 131:30]
  wire  dbRdReqArb_io_in_0_valid; // @[DCache.scala 137:28]
  wire [8:0] dbRdReqArb_io_in_0_bits_set; // @[DCache.scala 137:28]
  wire  dbRdReqArb_io_in_1_ready; // @[DCache.scala 137:28]
  wire  dbRdReqArb_io_in_1_valid; // @[DCache.scala 137:28]
  wire [8:0] dbRdReqArb_io_in_1_bits_set; // @[DCache.scala 137:28]
  wire  dbRdReqArb_io_out_valid; // @[DCache.scala 137:28]
  wire [8:0] dbRdReqArb_io_out_bits_set; // @[DCache.scala 137:28]
  wire  dirRdReqArb_io_in_0_valid; // @[DCache.scala 142:29]
  wire [31:0] dirRdReqArb_io_in_0_bits_addr; // @[DCache.scala 142:29]
  wire  dirRdReqArb_io_in_1_ready; // @[DCache.scala 142:29]
  wire  dirRdReqArb_io_in_1_valid; // @[DCache.scala 142:29]
  wire [31:0] dirRdReqArb_io_in_1_bits_addr; // @[DCache.scala 142:29]
  wire  dirRdReqArb_io_out_valid; // @[DCache.scala 142:29]
  wire [31:0] dirRdReqArb_io_out_bits_addr; // @[DCache.scala 142:29]
  wire  dataBankWrArb_io_in_0_valid; // @[DCache.scala 148:31]
  wire [8:0] dataBankWrArb_io_in_0_bits_set; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_0_bits_data_0; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_0_bits_data_1; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_0_bits_data_2; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_0_bits_data_3; // @[DCache.scala 148:31]
  wire [3:0] dataBankWrArb_io_in_0_bits_blockMask; // @[DCache.scala 148:31]
  wire [3:0] dataBankWrArb_io_in_0_bits_way; // @[DCache.scala 148:31]
  wire  dataBankWrArb_io_in_1_ready; // @[DCache.scala 148:31]
  wire  dataBankWrArb_io_in_1_valid; // @[DCache.scala 148:31]
  wire [8:0] dataBankWrArb_io_in_1_bits_set; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_1_bits_data_0; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_1_bits_data_1; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_1_bits_data_2; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_1_bits_data_3; // @[DCache.scala 148:31]
  wire [3:0] dataBankWrArb_io_in_1_bits_way; // @[DCache.scala 148:31]
  wire  dataBankWrArb_io_in_2_ready; // @[DCache.scala 148:31]
  wire  dataBankWrArb_io_in_2_valid; // @[DCache.scala 148:31]
  wire [8:0] dataBankWrArb_io_in_2_bits_set; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_2_bits_data_0; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_2_bits_data_1; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_2_bits_data_2; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_in_2_bits_data_3; // @[DCache.scala 148:31]
  wire [3:0] dataBankWrArb_io_in_2_bits_blockMask; // @[DCache.scala 148:31]
  wire [3:0] dataBankWrArb_io_in_2_bits_way; // @[DCache.scala 148:31]
  wire  dataBankWrArb_io_out_valid; // @[DCache.scala 148:31]
  wire [8:0] dataBankWrArb_io_out_bits_set; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_out_bits_data_0; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_out_bits_data_1; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_out_bits_data_2; // @[DCache.scala 148:31]
  wire [31:0] dataBankWrArb_io_out_bits_data_3; // @[DCache.scala 148:31]
  wire [3:0] dataBankWrArb_io_out_bits_blockMask; // @[DCache.scala 148:31]
  wire [3:0] dataBankWrArb_io_out_bits_way; // @[DCache.scala 148:31]
  wire  dirWrArb_io_in_0_valid; // @[DCache.scala 154:26]
  wire [31:0] dirWrArb_io_in_0_bits_addr; // @[DCache.scala 154:26]
  wire [3:0] dirWrArb_io_in_0_bits_way; // @[DCache.scala 154:26]
  wire  dirWrArb_io_in_1_ready; // @[DCache.scala 154:26]
  wire  dirWrArb_io_in_1_valid; // @[DCache.scala 154:26]
  wire [31:0] dirWrArb_io_in_1_bits_addr; // @[DCache.scala 154:26]
  wire [3:0] dirWrArb_io_in_1_bits_way; // @[DCache.scala 154:26]
  wire  dirWrArb_io_in_2_ready; // @[DCache.scala 154:26]
  wire  dirWrArb_io_in_2_valid; // @[DCache.scala 154:26]
  wire [31:0] dirWrArb_io_in_2_bits_addr; // @[DCache.scala 154:26]
  wire [3:0] dirWrArb_io_in_2_bits_way; // @[DCache.scala 154:26]
  wire  dirWrArb_io_out_valid; // @[DCache.scala 154:26]
  wire [31:0] dirWrArb_io_out_bits_addr; // @[DCache.scala 154:26]
  wire [3:0] dirWrArb_io_out_bits_way; // @[DCache.scala 154:26]
  wire [1:0] dirWrArb_io_out_bits_meta; // @[DCache.scala 154:26]
  LoadPipe loadPipe ( // @[DCache.scala 82:26]
    .clock(loadPipe_clock),
    .reset(loadPipe_reset),
    .io_load_req_ready(loadPipe_io_load_req_ready),
    .io_load_req_valid(loadPipe_io_load_req_valid),
    .io_load_req_bits_addr(loadPipe_io_load_req_bits_addr),
    .io_load_resp_ready(loadPipe_io_load_resp_ready),
    .io_load_resp_valid(loadPipe_io_load_resp_valid),
    .io_load_resp_bits_data(loadPipe_io_load_resp_bits_data),
    .io_dir_req_ready(loadPipe_io_dir_req_ready),
    .io_dir_req_valid(loadPipe_io_dir_req_valid),
    .io_dir_req_bits_addr(loadPipe_io_dir_req_bits_addr),
    .io_dir_resp_bits_hit(loadPipe_io_dir_resp_bits_hit),
    .io_dir_resp_bits_chosenWay(loadPipe_io_dir_resp_bits_chosenWay),
    .io_dir_resp_bits_isDirtyWay(loadPipe_io_dir_resp_bits_isDirtyWay),
    .io_dir_resp_bits_tagRdVec_0(loadPipe_io_dir_resp_bits_tagRdVec_0),
    .io_dir_resp_bits_tagRdVec_1(loadPipe_io_dir_resp_bits_tagRdVec_1),
    .io_dir_resp_bits_tagRdVec_2(loadPipe_io_dir_resp_bits_tagRdVec_2),
    .io_dir_resp_bits_tagRdVec_3(loadPipe_io_dir_resp_bits_tagRdVec_3),
    .io_dataBank_req_ready(loadPipe_io_dataBank_req_ready),
    .io_dataBank_req_valid(loadPipe_io_dataBank_req_valid),
    .io_dataBank_req_bits_set(loadPipe_io_dataBank_req_bits_set),
    .io_dataBank_resp_0_0(loadPipe_io_dataBank_resp_0_0),
    .io_dataBank_resp_0_1(loadPipe_io_dataBank_resp_0_1),
    .io_dataBank_resp_0_2(loadPipe_io_dataBank_resp_0_2),
    .io_dataBank_resp_0_3(loadPipe_io_dataBank_resp_0_3),
    .io_dataBank_resp_1_0(loadPipe_io_dataBank_resp_1_0),
    .io_dataBank_resp_1_1(loadPipe_io_dataBank_resp_1_1),
    .io_dataBank_resp_1_2(loadPipe_io_dataBank_resp_1_2),
    .io_dataBank_resp_1_3(loadPipe_io_dataBank_resp_1_3),
    .io_dataBank_resp_2_0(loadPipe_io_dataBank_resp_2_0),
    .io_dataBank_resp_2_1(loadPipe_io_dataBank_resp_2_1),
    .io_dataBank_resp_2_2(loadPipe_io_dataBank_resp_2_2),
    .io_dataBank_resp_2_3(loadPipe_io_dataBank_resp_2_3),
    .io_dataBank_resp_3_0(loadPipe_io_dataBank_resp_3_0),
    .io_dataBank_resp_3_1(loadPipe_io_dataBank_resp_3_1),
    .io_dataBank_resp_3_2(loadPipe_io_dataBank_resp_3_2),
    .io_dataBank_resp_3_3(loadPipe_io_dataBank_resp_3_3),
    .io_mshr_ready(loadPipe_io_mshr_ready),
    .io_mshr_valid(loadPipe_io_mshr_valid),
    .io_mshr_bits_addr(loadPipe_io_mshr_bits_addr),
    .io_mshr_bits_dirInfo_hit(loadPipe_io_mshr_bits_dirInfo_hit),
    .io_mshr_bits_dirInfo_chosenWay(loadPipe_io_mshr_bits_dirInfo_chosenWay),
    .io_mshr_bits_dirInfo_isDirtyWay(loadPipe_io_mshr_bits_dirInfo_isDirtyWay),
    .io_mshr_bits_dirtyTag(loadPipe_io_mshr_bits_dirtyTag),
    .io_mshr_bits_data_0(loadPipe_io_mshr_bits_data_0),
    .io_mshr_bits_data_1(loadPipe_io_mshr_bits_data_1),
    .io_mshr_bits_data_2(loadPipe_io_mshr_bits_data_2),
    .io_mshr_bits_data_3(loadPipe_io_mshr_bits_data_3)
  );
  StorePipe storePipe ( // @[DCache.scala 83:27]
    .clock(storePipe_clock),
    .reset(storePipe_reset),
    .io_store_req_ready(storePipe_io_store_req_ready),
    .io_store_req_valid(storePipe_io_store_req_valid),
    .io_store_req_bits_addr(storePipe_io_store_req_bits_addr),
    .io_store_req_bits_data(storePipe_io_store_req_bits_data),
    .io_store_req_bits_mask(storePipe_io_store_req_bits_mask),
    .io_store_resp_ready(storePipe_io_store_resp_ready),
    .io_store_resp_valid(storePipe_io_store_resp_valid),
    .io_dir_read_req_valid(storePipe_io_dir_read_req_valid),
    .io_dir_read_req_bits_addr(storePipe_io_dir_read_req_bits_addr),
    .io_dir_read_resp_bits_hit(storePipe_io_dir_read_resp_bits_hit),
    .io_dir_read_resp_bits_chosenWay(storePipe_io_dir_read_resp_bits_chosenWay),
    .io_dir_read_resp_bits_isDirtyWay(storePipe_io_dir_read_resp_bits_isDirtyWay),
    .io_dir_read_resp_bits_tagRdVec_0(storePipe_io_dir_read_resp_bits_tagRdVec_0),
    .io_dir_read_resp_bits_tagRdVec_1(storePipe_io_dir_read_resp_bits_tagRdVec_1),
    .io_dir_read_resp_bits_tagRdVec_2(storePipe_io_dir_read_resp_bits_tagRdVec_2),
    .io_dir_read_resp_bits_tagRdVec_3(storePipe_io_dir_read_resp_bits_tagRdVec_3),
    .io_dir_write_req_valid(storePipe_io_dir_write_req_valid),
    .io_dir_write_req_bits_addr(storePipe_io_dir_write_req_bits_addr),
    .io_dir_write_req_bits_way(storePipe_io_dir_write_req_bits_way),
    .io_dataBank_read_req_valid(storePipe_io_dataBank_read_req_valid),
    .io_dataBank_read_req_bits_set(storePipe_io_dataBank_read_req_bits_set),
    .io_dataBank_read_resp_0_0(storePipe_io_dataBank_read_resp_0_0),
    .io_dataBank_read_resp_0_1(storePipe_io_dataBank_read_resp_0_1),
    .io_dataBank_read_resp_0_2(storePipe_io_dataBank_read_resp_0_2),
    .io_dataBank_read_resp_0_3(storePipe_io_dataBank_read_resp_0_3),
    .io_dataBank_read_resp_1_0(storePipe_io_dataBank_read_resp_1_0),
    .io_dataBank_read_resp_1_1(storePipe_io_dataBank_read_resp_1_1),
    .io_dataBank_read_resp_1_2(storePipe_io_dataBank_read_resp_1_2),
    .io_dataBank_read_resp_1_3(storePipe_io_dataBank_read_resp_1_3),
    .io_dataBank_read_resp_2_0(storePipe_io_dataBank_read_resp_2_0),
    .io_dataBank_read_resp_2_1(storePipe_io_dataBank_read_resp_2_1),
    .io_dataBank_read_resp_2_2(storePipe_io_dataBank_read_resp_2_2),
    .io_dataBank_read_resp_2_3(storePipe_io_dataBank_read_resp_2_3),
    .io_dataBank_read_resp_3_0(storePipe_io_dataBank_read_resp_3_0),
    .io_dataBank_read_resp_3_1(storePipe_io_dataBank_read_resp_3_1),
    .io_dataBank_read_resp_3_2(storePipe_io_dataBank_read_resp_3_2),
    .io_dataBank_read_resp_3_3(storePipe_io_dataBank_read_resp_3_3),
    .io_dataBank_write_req_valid(storePipe_io_dataBank_write_req_valid),
    .io_dataBank_write_req_bits_set(storePipe_io_dataBank_write_req_bits_set),
    .io_dataBank_write_req_bits_data_0(storePipe_io_dataBank_write_req_bits_data_0),
    .io_dataBank_write_req_bits_data_1(storePipe_io_dataBank_write_req_bits_data_1),
    .io_dataBank_write_req_bits_data_2(storePipe_io_dataBank_write_req_bits_data_2),
    .io_dataBank_write_req_bits_data_3(storePipe_io_dataBank_write_req_bits_data_3),
    .io_dataBank_write_req_bits_blockMask(storePipe_io_dataBank_write_req_bits_blockMask),
    .io_dataBank_write_req_bits_way(storePipe_io_dataBank_write_req_bits_way),
    .io_mshr_ready(storePipe_io_mshr_ready),
    .io_mshr_valid(storePipe_io_mshr_valid),
    .io_mshr_bits_addr(storePipe_io_mshr_bits_addr),
    .io_mshr_bits_dirInfo_hit(storePipe_io_mshr_bits_dirInfo_hit),
    .io_mshr_bits_dirInfo_chosenWay(storePipe_io_mshr_bits_dirInfo_chosenWay),
    .io_mshr_bits_dirInfo_isDirtyWay(storePipe_io_mshr_bits_dirInfo_isDirtyWay),
    .io_mshr_bits_dirtyTag(storePipe_io_mshr_bits_dirtyTag),
    .io_mshr_bits_data_0(storePipe_io_mshr_bits_data_0),
    .io_mshr_bits_data_1(storePipe_io_mshr_bits_data_1),
    .io_mshr_bits_data_2(storePipe_io_mshr_bits_data_2),
    .io_mshr_bits_data_3(storePipe_io_mshr_bits_data_3),
    .io_mshr_bits_storeData(storePipe_io_mshr_bits_storeData),
    .io_mshr_bits_storeMask(storePipe_io_mshr_bits_storeMask),
    .io_flush(storePipe_io_flush)
  );
  MSHR mshr ( // @[DCache.scala 84:22]
    .clock(mshr_clock),
    .reset(mshr_reset),
    .io_req_ready(mshr_io_req_ready),
    .io_req_valid(mshr_io_req_valid),
    .io_req_bits_addr(mshr_io_req_bits_addr),
    .io_req_bits_dirInfo_hit(mshr_io_req_bits_dirInfo_hit),
    .io_req_bits_dirInfo_chosenWay(mshr_io_req_bits_dirInfo_chosenWay),
    .io_req_bits_dirInfo_isDirtyWay(mshr_io_req_bits_dirInfo_isDirtyWay),
    .io_req_bits_dirtyTag(mshr_io_req_bits_dirtyTag),
    .io_req_bits_data_0(mshr_io_req_bits_data_0),
    .io_req_bits_data_1(mshr_io_req_bits_data_1),
    .io_req_bits_data_2(mshr_io_req_bits_data_2),
    .io_req_bits_data_3(mshr_io_req_bits_data_3),
    .io_req_bits_isStore(mshr_io_req_bits_isStore),
    .io_req_bits_storeData(mshr_io_req_bits_storeData),
    .io_req_bits_storeMask(mshr_io_req_bits_storeMask),
    .io_resp_load_ready(mshr_io_resp_load_ready),
    .io_resp_load_valid(mshr_io_resp_load_valid),
    .io_resp_load_bits_data(mshr_io_resp_load_bits_data),
    .io_resp_store_ready(mshr_io_resp_store_ready),
    .io_resp_store_valid(mshr_io_resp_store_valid),
    .io_tasks_refill_req_valid(mshr_io_tasks_refill_req_valid),
    .io_tasks_refill_req_bits_addr(mshr_io_tasks_refill_req_bits_addr),
    .io_tasks_refill_req_bits_chosenWay(mshr_io_tasks_refill_req_bits_chosenWay),
    .io_tasks_refill_resp_ready(mshr_io_tasks_refill_resp_ready),
    .io_tasks_refill_resp_valid(mshr_io_tasks_refill_resp_valid),
    .io_tasks_refill_resp_bits_data(mshr_io_tasks_refill_resp_bits_data),
    .io_tasks_writeback_req_valid(mshr_io_tasks_writeback_req_valid),
    .io_tasks_writeback_req_bits_addr(mshr_io_tasks_writeback_req_bits_addr),
    .io_tasks_writeback_req_bits_dirtyTag(mshr_io_tasks_writeback_req_bits_dirtyTag),
    .io_tasks_writeback_req_bits_data_0(mshr_io_tasks_writeback_req_bits_data_0),
    .io_tasks_writeback_req_bits_data_1(mshr_io_tasks_writeback_req_bits_data_1),
    .io_tasks_writeback_req_bits_data_2(mshr_io_tasks_writeback_req_bits_data_2),
    .io_tasks_writeback_req_bits_data_3(mshr_io_tasks_writeback_req_bits_data_3),
    .io_tasks_writeback_resp_ready(mshr_io_tasks_writeback_resp_ready),
    .io_tasks_writeback_resp_valid(mshr_io_tasks_writeback_resp_valid),
    .io_dirWrite_req_ready(mshr_io_dirWrite_req_ready),
    .io_dirWrite_req_valid(mshr_io_dirWrite_req_valid),
    .io_dirWrite_req_bits_addr(mshr_io_dirWrite_req_bits_addr),
    .io_dirWrite_req_bits_way(mshr_io_dirWrite_req_bits_way),
    .io_dataWrite_req_ready(mshr_io_dataWrite_req_ready),
    .io_dataWrite_req_valid(mshr_io_dataWrite_req_valid),
    .io_dataWrite_req_bits_set(mshr_io_dataWrite_req_bits_set),
    .io_dataWrite_req_bits_data_0(mshr_io_dataWrite_req_bits_data_0),
    .io_dataWrite_req_bits_data_1(mshr_io_dataWrite_req_bits_data_1),
    .io_dataWrite_req_bits_data_2(mshr_io_dataWrite_req_bits_data_2),
    .io_dataWrite_req_bits_data_3(mshr_io_dataWrite_req_bits_data_3),
    .io_dataWrite_req_bits_blockMask(mshr_io_dataWrite_req_bits_blockMask),
    .io_dataWrite_req_bits_way(mshr_io_dataWrite_req_bits_way),
    .io_flush(mshr_io_flush)
  );
  RefillPipe_1 refillPipe ( // @[DCache.scala 85:28]
    .clock(refillPipe_clock),
    .reset(refillPipe_reset),
    .io_req_ready(refillPipe_io_req_ready),
    .io_req_valid(refillPipe_io_req_valid),
    .io_req_bits_addr(refillPipe_io_req_bits_addr),
    .io_req_bits_chosenWay(refillPipe_io_req_bits_chosenWay),
    .io_resp_valid(refillPipe_io_resp_valid),
    .io_resp_bits_data(refillPipe_io_resp_bits_data),
    .io_tlbus_req_ready(refillPipe_io_tlbus_req_ready),
    .io_tlbus_req_valid(refillPipe_io_tlbus_req_valid),
    .io_tlbus_req_bits_address(refillPipe_io_tlbus_req_bits_address),
    .io_tlbus_resp_ready(refillPipe_io_tlbus_resp_ready),
    .io_tlbus_resp_valid(refillPipe_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(refillPipe_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(refillPipe_io_tlbus_resp_bits_data),
    .io_dirWrite_req_ready(refillPipe_io_dirWrite_req_ready),
    .io_dirWrite_req_valid(refillPipe_io_dirWrite_req_valid),
    .io_dirWrite_req_bits_addr(refillPipe_io_dirWrite_req_bits_addr),
    .io_dirWrite_req_bits_way(refillPipe_io_dirWrite_req_bits_way),
    .io_dataWrite_req_ready(refillPipe_io_dataWrite_req_ready),
    .io_dataWrite_req_valid(refillPipe_io_dataWrite_req_valid),
    .io_dataWrite_req_bits_set(refillPipe_io_dataWrite_req_bits_set),
    .io_dataWrite_req_bits_data_0(refillPipe_io_dataWrite_req_bits_data_0),
    .io_dataWrite_req_bits_data_1(refillPipe_io_dataWrite_req_bits_data_1),
    .io_dataWrite_req_bits_data_2(refillPipe_io_dataWrite_req_bits_data_2),
    .io_dataWrite_req_bits_data_3(refillPipe_io_dataWrite_req_bits_data_3),
    .io_dataWrite_req_bits_way(refillPipe_io_dataWrite_req_bits_way)
  );
  WritebackQueue wb ( // @[DCache.scala 86:20]
    .clock(wb_clock),
    .reset(wb_reset),
    .io_req_ready(wb_io_req_ready),
    .io_req_valid(wb_io_req_valid),
    .io_req_bits_addr(wb_io_req_bits_addr),
    .io_req_bits_dirtyTag(wb_io_req_bits_dirtyTag),
    .io_req_bits_data_0(wb_io_req_bits_data_0),
    .io_req_bits_data_1(wb_io_req_bits_data_1),
    .io_req_bits_data_2(wb_io_req_bits_data_2),
    .io_req_bits_data_3(wb_io_req_bits_data_3),
    .io_resp_valid(wb_io_resp_valid),
    .io_tlbus_req_ready(wb_io_tlbus_req_ready),
    .io_tlbus_req_valid(wb_io_tlbus_req_valid),
    .io_tlbus_req_bits_address(wb_io_tlbus_req_bits_address),
    .io_tlbus_req_bits_data(wb_io_tlbus_req_bits_data),
    .io_tlbus_resp_ready(wb_io_tlbus_resp_ready),
    .io_tlbus_resp_valid(wb_io_tlbus_resp_valid)
  );
  DataBankArray_1 db ( // @[DCache.scala 87:20]
    .clock(db_clock),
    .reset(db_reset),
    .io_read_req_ready(db_io_read_req_ready),
    .io_read_req_valid(db_io_read_req_valid),
    .io_read_req_bits_set(db_io_read_req_bits_set),
    .io_read_resp_0_0(db_io_read_resp_0_0),
    .io_read_resp_0_1(db_io_read_resp_0_1),
    .io_read_resp_0_2(db_io_read_resp_0_2),
    .io_read_resp_0_3(db_io_read_resp_0_3),
    .io_read_resp_1_0(db_io_read_resp_1_0),
    .io_read_resp_1_1(db_io_read_resp_1_1),
    .io_read_resp_1_2(db_io_read_resp_1_2),
    .io_read_resp_1_3(db_io_read_resp_1_3),
    .io_read_resp_2_0(db_io_read_resp_2_0),
    .io_read_resp_2_1(db_io_read_resp_2_1),
    .io_read_resp_2_2(db_io_read_resp_2_2),
    .io_read_resp_2_3(db_io_read_resp_2_3),
    .io_read_resp_3_0(db_io_read_resp_3_0),
    .io_read_resp_3_1(db_io_read_resp_3_1),
    .io_read_resp_3_2(db_io_read_resp_3_2),
    .io_read_resp_3_3(db_io_read_resp_3_3),
    .io_write_req_ready(db_io_write_req_ready),
    .io_write_req_valid(db_io_write_req_valid),
    .io_write_req_bits_set(db_io_write_req_bits_set),
    .io_write_req_bits_data_0(db_io_write_req_bits_data_0),
    .io_write_req_bits_data_1(db_io_write_req_bits_data_1),
    .io_write_req_bits_data_2(db_io_write_req_bits_data_2),
    .io_write_req_bits_data_3(db_io_write_req_bits_data_3),
    .io_write_req_bits_blockMask(db_io_write_req_bits_blockMask),
    .io_write_req_bits_way(db_io_write_req_bits_way)
  );
  DCacheDirectory_1 dir ( // @[DCache.scala 88:21]
    .clock(dir_clock),
    .reset(dir_reset),
    .io_read_req_ready(dir_io_read_req_ready),
    .io_read_req_valid(dir_io_read_req_valid),
    .io_read_req_bits_addr(dir_io_read_req_bits_addr),
    .io_read_resp_bits_hit(dir_io_read_resp_bits_hit),
    .io_read_resp_bits_chosenWay(dir_io_read_resp_bits_chosenWay),
    .io_read_resp_bits_isDirtyWay(dir_io_read_resp_bits_isDirtyWay),
    .io_read_resp_bits_tagRdVec_0(dir_io_read_resp_bits_tagRdVec_0),
    .io_read_resp_bits_tagRdVec_1(dir_io_read_resp_bits_tagRdVec_1),
    .io_read_resp_bits_tagRdVec_2(dir_io_read_resp_bits_tagRdVec_2),
    .io_read_resp_bits_tagRdVec_3(dir_io_read_resp_bits_tagRdVec_3),
    .io_write_req_ready(dir_io_write_req_ready),
    .io_write_req_valid(dir_io_write_req_valid),
    .io_write_req_bits_addr(dir_io_write_req_bits_addr),
    .io_write_req_bits_way(dir_io_write_req_bits_way),
    .io_write_req_bits_meta(dir_io_write_req_bits_meta)
  );
  Arbiter_1 mshrReqArb ( // @[DCache.scala 109:28]
    .io_in_0_ready(mshrReqArb_io_in_0_ready),
    .io_in_0_valid(mshrReqArb_io_in_0_valid),
    .io_in_0_bits_addr(mshrReqArb_io_in_0_bits_addr),
    .io_in_0_bits_dirInfo_hit(mshrReqArb_io_in_0_bits_dirInfo_hit),
    .io_in_0_bits_dirInfo_chosenWay(mshrReqArb_io_in_0_bits_dirInfo_chosenWay),
    .io_in_0_bits_dirInfo_isDirtyWay(mshrReqArb_io_in_0_bits_dirInfo_isDirtyWay),
    .io_in_0_bits_dirtyTag(mshrReqArb_io_in_0_bits_dirtyTag),
    .io_in_0_bits_data_0(mshrReqArb_io_in_0_bits_data_0),
    .io_in_0_bits_data_1(mshrReqArb_io_in_0_bits_data_1),
    .io_in_0_bits_data_2(mshrReqArb_io_in_0_bits_data_2),
    .io_in_0_bits_data_3(mshrReqArb_io_in_0_bits_data_3),
    .io_in_1_ready(mshrReqArb_io_in_1_ready),
    .io_in_1_valid(mshrReqArb_io_in_1_valid),
    .io_in_1_bits_addr(mshrReqArb_io_in_1_bits_addr),
    .io_in_1_bits_dirInfo_hit(mshrReqArb_io_in_1_bits_dirInfo_hit),
    .io_in_1_bits_dirInfo_chosenWay(mshrReqArb_io_in_1_bits_dirInfo_chosenWay),
    .io_in_1_bits_dirInfo_isDirtyWay(mshrReqArb_io_in_1_bits_dirInfo_isDirtyWay),
    .io_in_1_bits_dirtyTag(mshrReqArb_io_in_1_bits_dirtyTag),
    .io_in_1_bits_data_0(mshrReqArb_io_in_1_bits_data_0),
    .io_in_1_bits_data_1(mshrReqArb_io_in_1_bits_data_1),
    .io_in_1_bits_data_2(mshrReqArb_io_in_1_bits_data_2),
    .io_in_1_bits_data_3(mshrReqArb_io_in_1_bits_data_3),
    .io_in_1_bits_storeData(mshrReqArb_io_in_1_bits_storeData),
    .io_in_1_bits_storeMask(mshrReqArb_io_in_1_bits_storeMask),
    .io_out_ready(mshrReqArb_io_out_ready),
    .io_out_valid(mshrReqArb_io_out_valid),
    .io_out_bits_addr(mshrReqArb_io_out_bits_addr),
    .io_out_bits_dirInfo_hit(mshrReqArb_io_out_bits_dirInfo_hit),
    .io_out_bits_dirInfo_chosenWay(mshrReqArb_io_out_bits_dirInfo_chosenWay),
    .io_out_bits_dirInfo_isDirtyWay(mshrReqArb_io_out_bits_dirInfo_isDirtyWay),
    .io_out_bits_dirtyTag(mshrReqArb_io_out_bits_dirtyTag),
    .io_out_bits_data_0(mshrReqArb_io_out_bits_data_0),
    .io_out_bits_data_1(mshrReqArb_io_out_bits_data_1),
    .io_out_bits_data_2(mshrReqArb_io_out_bits_data_2),
    .io_out_bits_data_3(mshrReqArb_io_out_bits_data_3),
    .io_out_bits_isStore(mshrReqArb_io_out_bits_isStore),
    .io_out_bits_storeData(mshrReqArb_io_out_bits_storeData),
    .io_out_bits_storeMask(mshrReqArb_io_out_bits_storeMask)
  );
  Arbiter_2 tlbusReqArb ( // @[DCache.scala 114:29]
    .io_in_0_ready(tlbusReqArb_io_in_0_ready),
    .io_in_0_valid(tlbusReqArb_io_in_0_valid),
    .io_in_0_bits_address(tlbusReqArb_io_in_0_bits_address),
    .io_in_0_bits_data(tlbusReqArb_io_in_0_bits_data),
    .io_in_1_ready(tlbusReqArb_io_in_1_ready),
    .io_in_1_valid(tlbusReqArb_io_in_1_valid),
    .io_in_1_bits_address(tlbusReqArb_io_in_1_bits_address),
    .io_out_ready(tlbusReqArb_io_out_ready),
    .io_out_valid(tlbusReqArb_io_out_valid),
    .io_out_bits_opcode(tlbusReqArb_io_out_bits_opcode),
    .io_out_bits_address(tlbusReqArb_io_out_bits_address),
    .io_out_bits_data(tlbusReqArb_io_out_bits_data)
  );
  Arbiter_3 loadRespArb ( // @[DCache.scala 126:29]
    .io_in_0_ready(loadRespArb_io_in_0_ready),
    .io_in_0_valid(loadRespArb_io_in_0_valid),
    .io_in_0_bits_data(loadRespArb_io_in_0_bits_data),
    .io_in_1_ready(loadRespArb_io_in_1_ready),
    .io_in_1_valid(loadRespArb_io_in_1_valid),
    .io_in_1_bits_data(loadRespArb_io_in_1_bits_data),
    .io_out_ready(loadRespArb_io_out_ready),
    .io_out_valid(loadRespArb_io_out_valid),
    .io_out_bits_data(loadRespArb_io_out_bits_data)
  );
  Arbiter_4 storeRespArb ( // @[DCache.scala 131:30]
    .io_in_0_ready(storeRespArb_io_in_0_ready),
    .io_in_0_valid(storeRespArb_io_in_0_valid),
    .io_in_1_ready(storeRespArb_io_in_1_ready),
    .io_in_1_valid(storeRespArb_io_in_1_valid),
    .io_out_ready(storeRespArb_io_out_ready),
    .io_out_valid(storeRespArb_io_out_valid)
  );
  Arbiter_5 dbRdReqArb ( // @[DCache.scala 137:28]
    .io_in_0_valid(dbRdReqArb_io_in_0_valid),
    .io_in_0_bits_set(dbRdReqArb_io_in_0_bits_set),
    .io_in_1_ready(dbRdReqArb_io_in_1_ready),
    .io_in_1_valid(dbRdReqArb_io_in_1_valid),
    .io_in_1_bits_set(dbRdReqArb_io_in_1_bits_set),
    .io_out_valid(dbRdReqArb_io_out_valid),
    .io_out_bits_set(dbRdReqArb_io_out_bits_set)
  );
  Arbiter_6 dirRdReqArb ( // @[DCache.scala 142:29]
    .io_in_0_valid(dirRdReqArb_io_in_0_valid),
    .io_in_0_bits_addr(dirRdReqArb_io_in_0_bits_addr),
    .io_in_1_ready(dirRdReqArb_io_in_1_ready),
    .io_in_1_valid(dirRdReqArb_io_in_1_valid),
    .io_in_1_bits_addr(dirRdReqArb_io_in_1_bits_addr),
    .io_out_valid(dirRdReqArb_io_out_valid),
    .io_out_bits_addr(dirRdReqArb_io_out_bits_addr)
  );
  Arbiter_7 dataBankWrArb ( // @[DCache.scala 148:31]
    .io_in_0_valid(dataBankWrArb_io_in_0_valid),
    .io_in_0_bits_set(dataBankWrArb_io_in_0_bits_set),
    .io_in_0_bits_data_0(dataBankWrArb_io_in_0_bits_data_0),
    .io_in_0_bits_data_1(dataBankWrArb_io_in_0_bits_data_1),
    .io_in_0_bits_data_2(dataBankWrArb_io_in_0_bits_data_2),
    .io_in_0_bits_data_3(dataBankWrArb_io_in_0_bits_data_3),
    .io_in_0_bits_blockMask(dataBankWrArb_io_in_0_bits_blockMask),
    .io_in_0_bits_way(dataBankWrArb_io_in_0_bits_way),
    .io_in_1_ready(dataBankWrArb_io_in_1_ready),
    .io_in_1_valid(dataBankWrArb_io_in_1_valid),
    .io_in_1_bits_set(dataBankWrArb_io_in_1_bits_set),
    .io_in_1_bits_data_0(dataBankWrArb_io_in_1_bits_data_0),
    .io_in_1_bits_data_1(dataBankWrArb_io_in_1_bits_data_1),
    .io_in_1_bits_data_2(dataBankWrArb_io_in_1_bits_data_2),
    .io_in_1_bits_data_3(dataBankWrArb_io_in_1_bits_data_3),
    .io_in_1_bits_way(dataBankWrArb_io_in_1_bits_way),
    .io_in_2_ready(dataBankWrArb_io_in_2_ready),
    .io_in_2_valid(dataBankWrArb_io_in_2_valid),
    .io_in_2_bits_set(dataBankWrArb_io_in_2_bits_set),
    .io_in_2_bits_data_0(dataBankWrArb_io_in_2_bits_data_0),
    .io_in_2_bits_data_1(dataBankWrArb_io_in_2_bits_data_1),
    .io_in_2_bits_data_2(dataBankWrArb_io_in_2_bits_data_2),
    .io_in_2_bits_data_3(dataBankWrArb_io_in_2_bits_data_3),
    .io_in_2_bits_blockMask(dataBankWrArb_io_in_2_bits_blockMask),
    .io_in_2_bits_way(dataBankWrArb_io_in_2_bits_way),
    .io_out_valid(dataBankWrArb_io_out_valid),
    .io_out_bits_set(dataBankWrArb_io_out_bits_set),
    .io_out_bits_data_0(dataBankWrArb_io_out_bits_data_0),
    .io_out_bits_data_1(dataBankWrArb_io_out_bits_data_1),
    .io_out_bits_data_2(dataBankWrArb_io_out_bits_data_2),
    .io_out_bits_data_3(dataBankWrArb_io_out_bits_data_3),
    .io_out_bits_blockMask(dataBankWrArb_io_out_bits_blockMask),
    .io_out_bits_way(dataBankWrArb_io_out_bits_way)
  );
  Arbiter_8 dirWrArb ( // @[DCache.scala 154:26]
    .io_in_0_valid(dirWrArb_io_in_0_valid),
    .io_in_0_bits_addr(dirWrArb_io_in_0_bits_addr),
    .io_in_0_bits_way(dirWrArb_io_in_0_bits_way),
    .io_in_1_ready(dirWrArb_io_in_1_ready),
    .io_in_1_valid(dirWrArb_io_in_1_valid),
    .io_in_1_bits_addr(dirWrArb_io_in_1_bits_addr),
    .io_in_1_bits_way(dirWrArb_io_in_1_bits_way),
    .io_in_2_ready(dirWrArb_io_in_2_ready),
    .io_in_2_valid(dirWrArb_io_in_2_valid),
    .io_in_2_bits_addr(dirWrArb_io_in_2_bits_addr),
    .io_in_2_bits_way(dirWrArb_io_in_2_bits_way),
    .io_out_valid(dirWrArb_io_out_valid),
    .io_out_bits_addr(dirWrArb_io_out_bits_addr),
    .io_out_bits_way(dirWrArb_io_out_bits_way),
    .io_out_bits_meta(dirWrArb_io_out_bits_meta)
  );
  assign io_read_req_ready = loadPipe_io_load_req_ready; // @[DCache.scala 101:26]
  assign io_read_resp_valid = loadRespArb_io_out_valid; // @[DCache.scala 129:18]
  assign io_read_resp_bits_data = loadRespArb_io_out_bits_data; // @[DCache.scala 129:18]
  assign io_write_req_ready = storePipe_io_store_req_ready; // @[DCache.scala 102:28]
  assign io_write_resp_valid = storeRespArb_io_out_valid; // @[DCache.scala 134:19]
  assign io_tlbus_req_valid = tlbusReqArb_io_out_valid; // @[DCache.scala 117:18]
  assign io_tlbus_req_bits_opcode = tlbusReqArb_io_out_bits_opcode; // @[DCache.scala 117:18]
  assign io_tlbus_req_bits_address = tlbusReqArb_io_out_bits_address; // @[DCache.scala 117:18]
  assign io_tlbus_req_bits_data = tlbusReqArb_io_out_bits_data; // @[DCache.scala 117:18]
  assign loadPipe_clock = clock;
  assign loadPipe_reset = reset;
  assign loadPipe_io_load_req_valid = io_read_req_valid; // @[DCache.scala 101:26]
  assign loadPipe_io_load_req_bits_addr = io_read_req_bits_addr; // @[DCache.scala 101:26]
  assign loadPipe_io_load_resp_ready = loadRespArb_io_in_0_ready; // @[DCache.scala 127:26]
  assign loadPipe_io_dir_req_ready = dirRdReqArb_io_in_1_ready; // @[DCache.scala 144:26]
  assign loadPipe_io_dir_resp_bits_hit = dir_io_read_resp_bits_hit; // @[DCache.scala 94:31]
  assign loadPipe_io_dir_resp_bits_chosenWay = dir_io_read_resp_bits_chosenWay; // @[DCache.scala 94:31]
  assign loadPipe_io_dir_resp_bits_isDirtyWay = dir_io_read_resp_bits_isDirtyWay; // @[DCache.scala 94:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_0 = dir_io_read_resp_bits_tagRdVec_0; // @[DCache.scala 94:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_1 = dir_io_read_resp_bits_tagRdVec_1; // @[DCache.scala 94:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_2 = dir_io_read_resp_bits_tagRdVec_2; // @[DCache.scala 94:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_3 = dir_io_read_resp_bits_tagRdVec_3; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_req_ready = dbRdReqArb_io_in_1_ready; // @[DCache.scala 139:25]
  assign loadPipe_io_dataBank_resp_0_0 = db_io_read_resp_0_0; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_0_1 = db_io_read_resp_0_1; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_0_2 = db_io_read_resp_0_2; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_0_3 = db_io_read_resp_0_3; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_1_0 = db_io_read_resp_1_0; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_1_1 = db_io_read_resp_1_1; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_1_2 = db_io_read_resp_1_2; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_1_3 = db_io_read_resp_1_3; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_2_0 = db_io_read_resp_2_0; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_2_1 = db_io_read_resp_2_1; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_2_2 = db_io_read_resp_2_2; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_2_3 = db_io_read_resp_2_3; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_3_0 = db_io_read_resp_3_0; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_3_1 = db_io_read_resp_3_1; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_3_2 = db_io_read_resp_3_2; // @[DCache.scala 98:31]
  assign loadPipe_io_dataBank_resp_3_3 = db_io_read_resp_3_3; // @[DCache.scala 98:31]
  assign loadPipe_io_mshr_ready = mshrReqArb_io_in_0_ready; // @[DCache.scala 110:25]
  assign storePipe_clock = clock;
  assign storePipe_reset = reset;
  assign storePipe_io_store_req_valid = io_write_req_valid; // @[DCache.scala 102:28]
  assign storePipe_io_store_req_bits_addr = io_write_req_bits_addr; // @[DCache.scala 102:28]
  assign storePipe_io_store_req_bits_data = io_write_req_bits_data; // @[DCache.scala 102:28]
  assign storePipe_io_store_req_bits_mask = io_write_req_bits_mask; // @[DCache.scala 102:28]
  assign storePipe_io_store_resp_ready = storeRespArb_io_in_0_ready; // @[DCache.scala 132:27]
  assign storePipe_io_dir_read_resp_bits_hit = dir_io_read_resp_bits_hit; // @[DCache.scala 96:37]
  assign storePipe_io_dir_read_resp_bits_chosenWay = dir_io_read_resp_bits_chosenWay; // @[DCache.scala 96:37]
  assign storePipe_io_dir_read_resp_bits_isDirtyWay = dir_io_read_resp_bits_isDirtyWay; // @[DCache.scala 96:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_0 = dir_io_read_resp_bits_tagRdVec_0; // @[DCache.scala 96:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_1 = dir_io_read_resp_bits_tagRdVec_1; // @[DCache.scala 96:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_2 = dir_io_read_resp_bits_tagRdVec_2; // @[DCache.scala 96:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_3 = dir_io_read_resp_bits_tagRdVec_3; // @[DCache.scala 96:37]
  assign storePipe_io_dataBank_read_resp_0_0 = db_io_read_resp_0_0; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_0_1 = db_io_read_resp_0_1; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_0_2 = db_io_read_resp_0_2; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_0_3 = db_io_read_resp_0_3; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_1_0 = db_io_read_resp_1_0; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_1_1 = db_io_read_resp_1_1; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_1_2 = db_io_read_resp_1_2; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_1_3 = db_io_read_resp_1_3; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_2_0 = db_io_read_resp_2_0; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_2_1 = db_io_read_resp_2_1; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_2_2 = db_io_read_resp_2_2; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_2_3 = db_io_read_resp_2_3; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_3_0 = db_io_read_resp_3_0; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_3_1 = db_io_read_resp_3_1; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_3_2 = db_io_read_resp_3_2; // @[DCache.scala 99:37]
  assign storePipe_io_dataBank_read_resp_3_3 = db_io_read_resp_3_3; // @[DCache.scala 99:37]
  assign storePipe_io_mshr_ready = mshrReqArb_io_in_1_ready; // @[DCache.scala 111:25]
  assign storePipe_io_flush = io_flush; // @[DCache.scala 90:24]
  assign mshr_clock = clock;
  assign mshr_reset = reset;
  assign mshr_io_req_valid = mshrReqArb_io_out_valid; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_addr = mshrReqArb_io_out_bits_addr; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_dirInfo_hit = mshrReqArb_io_out_bits_dirInfo_hit; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_dirInfo_chosenWay = mshrReqArb_io_out_bits_dirInfo_chosenWay; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_dirInfo_isDirtyWay = mshrReqArb_io_out_bits_dirInfo_isDirtyWay; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_dirtyTag = mshrReqArb_io_out_bits_dirtyTag; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_data_0 = mshrReqArb_io_out_bits_data_0; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_data_1 = mshrReqArb_io_out_bits_data_1; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_data_2 = mshrReqArb_io_out_bits_data_2; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_data_3 = mshrReqArb_io_out_bits_data_3; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_isStore = mshrReqArb_io_out_bits_isStore; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_storeData = mshrReqArb_io_out_bits_storeData; // @[DCache.scala 112:17]
  assign mshr_io_req_bits_storeMask = mshrReqArb_io_out_bits_storeMask; // @[DCache.scala 112:17]
  assign mshr_io_resp_load_ready = loadRespArb_io_in_1_ready; // @[DCache.scala 128:26]
  assign mshr_io_resp_store_ready = storeRespArb_io_in_1_ready; // @[DCache.scala 133:27]
  assign mshr_io_tasks_refill_resp_valid = refillPipe_io_resp_valid; // @[DCache.scala 105:31]
  assign mshr_io_tasks_refill_resp_bits_data = refillPipe_io_resp_bits_data; // @[DCache.scala 105:31]
  assign mshr_io_tasks_writeback_resp_valid = wb_io_resp_valid; // @[DCache.scala 107:34]
  assign mshr_io_dirWrite_req_ready = dirWrArb_io_in_2_ready; // @[DCache.scala 157:23]
  assign mshr_io_dataWrite_req_ready = dataBankWrArb_io_in_2_ready; // @[DCache.scala 151:28]
  assign mshr_io_flush = io_flush; // @[DCache.scala 91:19]
  assign refillPipe_clock = clock;
  assign refillPipe_reset = reset;
  assign refillPipe_io_req_valid = mshr_io_tasks_refill_req_valid; // @[DCache.scala 104:30]
  assign refillPipe_io_req_bits_addr = mshr_io_tasks_refill_req_bits_addr; // @[DCache.scala 104:30]
  assign refillPipe_io_req_bits_chosenWay = mshr_io_tasks_refill_req_bits_chosenWay; // @[DCache.scala 104:30]
  assign refillPipe_io_tlbus_req_ready = tlbusReqArb_io_in_1_ready; // @[DCache.scala 116:26]
  assign refillPipe_io_tlbus_resp_valid = io_tlbus_resp_valid; // @[DCache.scala 121:36]
  assign refillPipe_io_tlbus_resp_bits_opcode = io_tlbus_resp_bits_opcode; // @[DCache.scala 122:35]
  assign refillPipe_io_tlbus_resp_bits_data = io_tlbus_resp_bits_data; // @[DCache.scala 122:35]
  assign refillPipe_io_dirWrite_req_ready = dirWrArb_io_in_1_ready; // @[DCache.scala 156:23]
  assign refillPipe_io_dataWrite_req_ready = dataBankWrArb_io_in_1_ready; // @[DCache.scala 150:28]
  assign wb_clock = clock;
  assign wb_reset = reset;
  assign wb_io_req_valid = mshr_io_tasks_writeback_req_valid; // @[DCache.scala 106:33]
  assign wb_io_req_bits_addr = mshr_io_tasks_writeback_req_bits_addr; // @[DCache.scala 106:33]
  assign wb_io_req_bits_dirtyTag = mshr_io_tasks_writeback_req_bits_dirtyTag; // @[DCache.scala 106:33]
  assign wb_io_req_bits_data_0 = mshr_io_tasks_writeback_req_bits_data_0; // @[DCache.scala 106:33]
  assign wb_io_req_bits_data_1 = mshr_io_tasks_writeback_req_bits_data_1; // @[DCache.scala 106:33]
  assign wb_io_req_bits_data_2 = mshr_io_tasks_writeback_req_bits_data_2; // @[DCache.scala 106:33]
  assign wb_io_req_bits_data_3 = mshr_io_tasks_writeback_req_bits_data_3; // @[DCache.scala 106:33]
  assign wb_io_tlbus_req_ready = tlbusReqArb_io_in_0_ready; // @[DCache.scala 115:26]
  assign wb_io_tlbus_resp_valid = io_tlbus_resp_valid; // @[DCache.scala 119:28]
  assign db_clock = clock;
  assign db_reset = reset;
  assign db_io_read_req_valid = dbRdReqArb_io_out_valid; // @[DCache.scala 140:20]
  assign db_io_read_req_bits_set = dbRdReqArb_io_out_bits_set; // @[DCache.scala 140:20]
  assign db_io_write_req_valid = dataBankWrArb_io_out_valid; // @[DCache.scala 152:21]
  assign db_io_write_req_bits_set = dataBankWrArb_io_out_bits_set; // @[DCache.scala 152:21]
  assign db_io_write_req_bits_data_0 = dataBankWrArb_io_out_bits_data_0; // @[DCache.scala 152:21]
  assign db_io_write_req_bits_data_1 = dataBankWrArb_io_out_bits_data_1; // @[DCache.scala 152:21]
  assign db_io_write_req_bits_data_2 = dataBankWrArb_io_out_bits_data_2; // @[DCache.scala 152:21]
  assign db_io_write_req_bits_data_3 = dataBankWrArb_io_out_bits_data_3; // @[DCache.scala 152:21]
  assign db_io_write_req_bits_blockMask = dataBankWrArb_io_out_bits_blockMask; // @[DCache.scala 152:21]
  assign db_io_write_req_bits_way = dataBankWrArb_io_out_bits_way; // @[DCache.scala 152:21]
  assign dir_clock = clock;
  assign dir_reset = reset;
  assign dir_io_read_req_valid = dirRdReqArb_io_out_valid; // @[DCache.scala 145:21]
  assign dir_io_read_req_bits_addr = dirRdReqArb_io_out_bits_addr; // @[DCache.scala 145:21]
  assign dir_io_write_req_valid = dirWrArb_io_out_valid; // @[DCache.scala 158:22]
  assign dir_io_write_req_bits_addr = dirWrArb_io_out_bits_addr; // @[DCache.scala 158:22]
  assign dir_io_write_req_bits_way = dirWrArb_io_out_bits_way; // @[DCache.scala 158:22]
  assign dir_io_write_req_bits_meta = dirWrArb_io_out_bits_meta; // @[DCache.scala 158:22]
  assign mshrReqArb_io_in_0_valid = loadPipe_io_mshr_valid; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_0_bits_addr = loadPipe_io_mshr_bits_addr; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_0_bits_dirInfo_hit = loadPipe_io_mshr_bits_dirInfo_hit; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_0_bits_dirInfo_chosenWay = loadPipe_io_mshr_bits_dirInfo_chosenWay; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_0_bits_dirInfo_isDirtyWay = loadPipe_io_mshr_bits_dirInfo_isDirtyWay; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_0_bits_dirtyTag = loadPipe_io_mshr_bits_dirtyTag; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_0_bits_data_0 = loadPipe_io_mshr_bits_data_0; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_0_bits_data_1 = loadPipe_io_mshr_bits_data_1; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_0_bits_data_2 = loadPipe_io_mshr_bits_data_2; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_0_bits_data_3 = loadPipe_io_mshr_bits_data_3; // @[DCache.scala 110:25]
  assign mshrReqArb_io_in_1_valid = storePipe_io_mshr_valid; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_addr = storePipe_io_mshr_bits_addr; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_dirInfo_hit = storePipe_io_mshr_bits_dirInfo_hit; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_dirInfo_chosenWay = storePipe_io_mshr_bits_dirInfo_chosenWay; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_dirInfo_isDirtyWay = storePipe_io_mshr_bits_dirInfo_isDirtyWay; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_dirtyTag = storePipe_io_mshr_bits_dirtyTag; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_data_0 = storePipe_io_mshr_bits_data_0; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_data_1 = storePipe_io_mshr_bits_data_1; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_data_2 = storePipe_io_mshr_bits_data_2; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_data_3 = storePipe_io_mshr_bits_data_3; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_storeData = storePipe_io_mshr_bits_storeData; // @[DCache.scala 111:25]
  assign mshrReqArb_io_in_1_bits_storeMask = storePipe_io_mshr_bits_storeMask; // @[DCache.scala 111:25]
  assign mshrReqArb_io_out_ready = mshr_io_req_ready; // @[DCache.scala 112:17]
  assign tlbusReqArb_io_in_0_valid = wb_io_tlbus_req_valid; // @[DCache.scala 115:26]
  assign tlbusReqArb_io_in_0_bits_address = wb_io_tlbus_req_bits_address; // @[DCache.scala 115:26]
  assign tlbusReqArb_io_in_0_bits_data = wb_io_tlbus_req_bits_data; // @[DCache.scala 115:26]
  assign tlbusReqArb_io_in_1_valid = refillPipe_io_tlbus_req_valid; // @[DCache.scala 116:26]
  assign tlbusReqArb_io_in_1_bits_address = refillPipe_io_tlbus_req_bits_address; // @[DCache.scala 116:26]
  assign tlbusReqArb_io_out_ready = io_tlbus_req_ready; // @[DCache.scala 117:18]
  assign loadRespArb_io_in_0_valid = loadPipe_io_load_resp_valid; // @[DCache.scala 127:26]
  assign loadRespArb_io_in_0_bits_data = loadPipe_io_load_resp_bits_data; // @[DCache.scala 127:26]
  assign loadRespArb_io_in_1_valid = mshr_io_resp_load_valid; // @[DCache.scala 128:26]
  assign loadRespArb_io_in_1_bits_data = mshr_io_resp_load_bits_data; // @[DCache.scala 128:26]
  assign loadRespArb_io_out_ready = io_read_resp_ready; // @[DCache.scala 129:18]
  assign storeRespArb_io_in_0_valid = storePipe_io_store_resp_valid; // @[DCache.scala 132:27]
  assign storeRespArb_io_in_1_valid = mshr_io_resp_store_valid; // @[DCache.scala 133:27]
  assign storeRespArb_io_out_ready = io_write_resp_ready; // @[DCache.scala 134:19]
  assign dbRdReqArb_io_in_0_valid = storePipe_io_dataBank_read_req_valid; // @[DCache.scala 138:25]
  assign dbRdReqArb_io_in_0_bits_set = storePipe_io_dataBank_read_req_bits_set; // @[DCache.scala 138:25]
  assign dbRdReqArb_io_in_1_valid = loadPipe_io_dataBank_req_valid; // @[DCache.scala 139:25]
  assign dbRdReqArb_io_in_1_bits_set = loadPipe_io_dataBank_req_bits_set; // @[DCache.scala 139:25]
  assign dirRdReqArb_io_in_0_valid = storePipe_io_dir_read_req_valid; // @[DCache.scala 143:26]
  assign dirRdReqArb_io_in_0_bits_addr = storePipe_io_dir_read_req_bits_addr; // @[DCache.scala 143:26]
  assign dirRdReqArb_io_in_1_valid = loadPipe_io_dir_req_valid; // @[DCache.scala 144:26]
  assign dirRdReqArb_io_in_1_bits_addr = loadPipe_io_dir_req_bits_addr; // @[DCache.scala 144:26]
  assign dataBankWrArb_io_in_0_valid = storePipe_io_dataBank_write_req_valid; // @[DCache.scala 149:28]
  assign dataBankWrArb_io_in_0_bits_set = storePipe_io_dataBank_write_req_bits_set; // @[DCache.scala 149:28]
  assign dataBankWrArb_io_in_0_bits_data_0 = storePipe_io_dataBank_write_req_bits_data_0; // @[DCache.scala 149:28]
  assign dataBankWrArb_io_in_0_bits_data_1 = storePipe_io_dataBank_write_req_bits_data_1; // @[DCache.scala 149:28]
  assign dataBankWrArb_io_in_0_bits_data_2 = storePipe_io_dataBank_write_req_bits_data_2; // @[DCache.scala 149:28]
  assign dataBankWrArb_io_in_0_bits_data_3 = storePipe_io_dataBank_write_req_bits_data_3; // @[DCache.scala 149:28]
  assign dataBankWrArb_io_in_0_bits_blockMask = storePipe_io_dataBank_write_req_bits_blockMask; // @[DCache.scala 149:28]
  assign dataBankWrArb_io_in_0_bits_way = storePipe_io_dataBank_write_req_bits_way; // @[DCache.scala 149:28]
  assign dataBankWrArb_io_in_1_valid = refillPipe_io_dataWrite_req_valid; // @[DCache.scala 150:28]
  assign dataBankWrArb_io_in_1_bits_set = refillPipe_io_dataWrite_req_bits_set; // @[DCache.scala 150:28]
  assign dataBankWrArb_io_in_1_bits_data_0 = refillPipe_io_dataWrite_req_bits_data_0; // @[DCache.scala 150:28]
  assign dataBankWrArb_io_in_1_bits_data_1 = refillPipe_io_dataWrite_req_bits_data_1; // @[DCache.scala 150:28]
  assign dataBankWrArb_io_in_1_bits_data_2 = refillPipe_io_dataWrite_req_bits_data_2; // @[DCache.scala 150:28]
  assign dataBankWrArb_io_in_1_bits_data_3 = refillPipe_io_dataWrite_req_bits_data_3; // @[DCache.scala 150:28]
  assign dataBankWrArb_io_in_1_bits_way = refillPipe_io_dataWrite_req_bits_way; // @[DCache.scala 150:28]
  assign dataBankWrArb_io_in_2_valid = mshr_io_dataWrite_req_valid; // @[DCache.scala 151:28]
  assign dataBankWrArb_io_in_2_bits_set = mshr_io_dataWrite_req_bits_set; // @[DCache.scala 151:28]
  assign dataBankWrArb_io_in_2_bits_data_0 = mshr_io_dataWrite_req_bits_data_0; // @[DCache.scala 151:28]
  assign dataBankWrArb_io_in_2_bits_data_1 = mshr_io_dataWrite_req_bits_data_1; // @[DCache.scala 151:28]
  assign dataBankWrArb_io_in_2_bits_data_2 = mshr_io_dataWrite_req_bits_data_2; // @[DCache.scala 151:28]
  assign dataBankWrArb_io_in_2_bits_data_3 = mshr_io_dataWrite_req_bits_data_3; // @[DCache.scala 151:28]
  assign dataBankWrArb_io_in_2_bits_blockMask = mshr_io_dataWrite_req_bits_blockMask; // @[DCache.scala 151:28]
  assign dataBankWrArb_io_in_2_bits_way = mshr_io_dataWrite_req_bits_way; // @[DCache.scala 151:28]
  assign dirWrArb_io_in_0_valid = storePipe_io_dir_write_req_valid; // @[DCache.scala 155:23]
  assign dirWrArb_io_in_0_bits_addr = storePipe_io_dir_write_req_bits_addr; // @[DCache.scala 155:23]
  assign dirWrArb_io_in_0_bits_way = storePipe_io_dir_write_req_bits_way; // @[DCache.scala 155:23]
  assign dirWrArb_io_in_1_valid = refillPipe_io_dirWrite_req_valid; // @[DCache.scala 156:23]
  assign dirWrArb_io_in_1_bits_addr = refillPipe_io_dirWrite_req_bits_addr; // @[DCache.scala 156:23]
  assign dirWrArb_io_in_1_bits_way = refillPipe_io_dirWrite_req_bits_way; // @[DCache.scala 156:23]
  assign dirWrArb_io_in_2_valid = mshr_io_dirWrite_req_valid; // @[DCache.scala 157:23]
  assign dirWrArb_io_in_2_bits_addr = mshr_io_dirWrite_req_bits_addr; // @[DCache.scala 157:23]
  assign dirWrArb_io_in_2_bits_way = mshr_io_dirWrite_req_bits_way; // @[DCache.scala 157:23]
endmodule
module TLBusArbiter(
  input        clock,
  input        reset,
  input        io_reqs_1,
  output [1:0] io_grantOH
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] owner; // @[Bus.scala 162:24]
  wire [3:0] _io_grantOH_T = 4'h1 << owner; // @[OneHot.scala 57:35]
  assign io_grantOH = _io_grantOH_T[1:0]; // @[Bus.scala 190:16]
  always @(posedge clock) begin
    if (reset) begin // @[Bus.scala 162:24]
      owner <= 2'h0; // @[Bus.scala 162:24]
    end else if (io_reqs_1) begin // @[Mux.scala 27:73]
      owner <= 2'h1;
    end else begin
      owner <= 2'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  owner = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBusMux(
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [31:0]  io_in_0_bits_address,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [2:0]   io_in_1_bits_opcode,
  input  [31:0]  io_in_1_bits_address,
  input  [127:0] io_in_1_bits_data,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_opcode,
  output [127:0] io_out_bits_size,
  output         io_out_bits_source,
  output [31:0]  io_out_bits_address,
  output [127:0] io_out_bits_data,
  input          io_choseOH_0,
  input          io_choseOH_1
);
  wire [31:0] _io_out_bits_T_9 = io_choseOH_0 ? io_in_0_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_bits_T_10 = io_choseOH_1 ? io_in_1_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [127:0] _io_out_bits_T_15 = io_choseOH_0 ? 128'h20 : 128'h0; // @[Mux.scala 27:73]
  wire [127:0] _io_out_bits_T_16 = io_choseOH_1 ? 128'h10 : 128'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_21 = io_choseOH_0 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_22 = io_choseOH_1 ? io_in_1_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  assign io_in_0_ready = io_out_ready & io_choseOH_0; // @[Bus.scala 132:80]
  assign io_in_1_ready = io_out_ready & io_choseOH_1; // @[Bus.scala 132:80]
  assign io_out_valid = io_choseOH_0 & io_in_0_valid | io_choseOH_1 & io_in_1_valid; // @[Mux.scala 27:73]
  assign io_out_bits_opcode = _io_out_bits_T_21 | _io_out_bits_T_22; // @[Mux.scala 27:73]
  assign io_out_bits_size = _io_out_bits_T_15 | _io_out_bits_T_16; // @[Mux.scala 27:73]
  assign io_out_bits_source = io_choseOH_1; // @[Mux.scala 27:73]
  assign io_out_bits_address = _io_out_bits_T_9 | _io_out_bits_T_10; // @[Mux.scala 27:73]
  assign io_out_bits_data = io_choseOH_1 ? io_in_1_bits_data : 128'h0; // @[Mux.scala 27:73]
endmodule
module Queue_6(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [2:0]   io_enq_bits_opcode,
  input  [127:0] io_enq_bits_size,
  input          io_enq_bits_source,
  input  [31:0]  io_enq_bits_address,
  input  [127:0] io_enq_bits_data,
  input          io_deq_ready,
  output         io_deq_valid,
  output [2:0]   io_deq_bits_opcode,
  output [127:0] io_deq_bits_size,
  output         io_deq_bits_source,
  output [31:0]  io_deq_bits_address,
  output [127:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_opcode_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 273:95]
  reg [127:0] ram_size [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [127:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [127:0] ram_size_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_source [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg [31:0] ram_address [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_address_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 273:95]
  reg [127:0] ram_data [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [127:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [127:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire  _GEN_19 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_19 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = enq_ptr_value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_opcode = empty ? io_enq_bits_opcode : ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_source = empty ? io_enq_bits_source : ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_address = empty ? io_enq_bits_address : ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[127:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_address[initvar] = _RAND_3[31:0];
  _RAND_4 = {4{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_data[initvar] = _RAND_4[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enq_ptr_value = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  deq_ptr_value = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLAddrDecode(
  input  [31:0] io_addr,
  output        io_choseOH_0,
  output        io_choseOH_1
);
  wire  valid = io_addr < 32'h10000000; // @[Bus.scala 201:42]
  wire  valid_1 = io_addr >= 32'h10000000 & io_addr < 32'h20000000; // @[Bus.scala 201:31]
  wire  _GEN_2 = valid_1 ? 1'h0 : 1'h1; // @[Bus.scala 211:68 212:20 214:20]
  assign io_choseOH_0 = valid | _GEN_2; // @[Bus.scala 209:62 210:20]
  assign io_choseOH_1 = valid ? 1'h0 : valid_1; // @[Bus.scala 209:62 210:20]
endmodule
module TLBusMux_1(
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [2:0]   io_in_0_bits_opcode,
  input  [127:0] io_in_0_bits_data,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_opcode,
  output [127:0] io_out_bits_data,
  input          io_choseOH_0
);
  assign io_in_0_ready = io_out_ready & io_choseOH_0; // @[Bus.scala 132:80]
  assign io_out_valid = io_choseOH_0 & io_in_0_valid; // @[Mux.scala 27:73]
  assign io_out_bits_opcode = io_choseOH_0 ? io_in_0_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  assign io_out_bits_data = io_choseOH_0 ? io_in_0_bits_data : 128'h0; // @[Mux.scala 27:73]
endmodule
module TLXbar(
  input          clock,
  input          reset,
  output         io_masterFace_in_0_ready,
  input          io_masterFace_in_0_valid,
  input  [31:0]  io_masterFace_in_0_bits_address,
  output         io_masterFace_in_1_ready,
  input          io_masterFace_in_1_valid,
  input  [2:0]   io_masterFace_in_1_bits_opcode,
  input  [31:0]  io_masterFace_in_1_bits_address,
  input  [127:0] io_masterFace_in_1_bits_data,
  output         io_masterFace_out_0_valid,
  output [2:0]   io_masterFace_out_0_bits_opcode,
  output [127:0] io_masterFace_out_0_bits_data,
  output         io_masterFace_out_1_valid,
  output [2:0]   io_masterFace_out_1_bits_opcode,
  output [127:0] io_masterFace_out_1_bits_data,
  input          io_slaveFace_in_0_ready,
  output         io_slaveFace_in_0_valid,
  output [2:0]   io_slaveFace_in_0_bits_opcode,
  output [127:0] io_slaveFace_in_0_bits_size,
  output [31:0]  io_slaveFace_in_0_bits_address,
  output [127:0] io_slaveFace_in_0_bits_data,
  output         io_slaveFace_out_0_ready,
  input          io_slaveFace_out_0_valid,
  input  [2:0]   io_slaveFace_out_0_bits_opcode,
  input  [127:0] io_slaveFace_out_0_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  reqArb_clock; // @[Bus.scala 233:24]
  wire  reqArb_reset; // @[Bus.scala 233:24]
  wire  reqArb_io_reqs_1; // @[Bus.scala 233:24]
  wire [1:0] reqArb_io_grantOH; // @[Bus.scala 233:24]
  wire  reqMux_io_in_0_ready; // @[Bus.scala 236:24]
  wire  reqMux_io_in_0_valid; // @[Bus.scala 236:24]
  wire [31:0] reqMux_io_in_0_bits_address; // @[Bus.scala 236:24]
  wire  reqMux_io_in_1_ready; // @[Bus.scala 236:24]
  wire  reqMux_io_in_1_valid; // @[Bus.scala 236:24]
  wire [2:0] reqMux_io_in_1_bits_opcode; // @[Bus.scala 236:24]
  wire [31:0] reqMux_io_in_1_bits_address; // @[Bus.scala 236:24]
  wire [127:0] reqMux_io_in_1_bits_data; // @[Bus.scala 236:24]
  wire  reqMux_io_out_ready; // @[Bus.scala 236:24]
  wire  reqMux_io_out_valid; // @[Bus.scala 236:24]
  wire [2:0] reqMux_io_out_bits_opcode; // @[Bus.scala 236:24]
  wire [127:0] reqMux_io_out_bits_size; // @[Bus.scala 236:24]
  wire  reqMux_io_out_bits_source; // @[Bus.scala 236:24]
  wire [31:0] reqMux_io_out_bits_address; // @[Bus.scala 236:24]
  wire [127:0] reqMux_io_out_bits_data; // @[Bus.scala 236:24]
  wire  reqMux_io_choseOH_0; // @[Bus.scala 236:24]
  wire  reqMux_io_choseOH_1; // @[Bus.scala 236:24]
  wire  buf__clock; // @[Bus.scala 242:21]
  wire  buf__reset; // @[Bus.scala 242:21]
  wire  buf__io_enq_ready; // @[Bus.scala 242:21]
  wire  buf__io_enq_valid; // @[Bus.scala 242:21]
  wire [2:0] buf__io_enq_bits_opcode; // @[Bus.scala 242:21]
  wire [127:0] buf__io_enq_bits_size; // @[Bus.scala 242:21]
  wire  buf__io_enq_bits_source; // @[Bus.scala 242:21]
  wire [31:0] buf__io_enq_bits_address; // @[Bus.scala 242:21]
  wire [127:0] buf__io_enq_bits_data; // @[Bus.scala 242:21]
  wire  buf__io_deq_ready; // @[Bus.scala 242:21]
  wire  buf__io_deq_valid; // @[Bus.scala 242:21]
  wire [2:0] buf__io_deq_bits_opcode; // @[Bus.scala 242:21]
  wire [127:0] buf__io_deq_bits_size; // @[Bus.scala 242:21]
  wire  buf__io_deq_bits_source; // @[Bus.scala 242:21]
  wire [31:0] buf__io_deq_bits_address; // @[Bus.scala 242:21]
  wire [127:0] buf__io_deq_bits_data; // @[Bus.scala 242:21]
  wire [31:0] addrDec_io_addr; // @[Bus.scala 265:25]
  wire  addrDec_io_choseOH_0; // @[Bus.scala 265:25]
  wire  addrDec_io_choseOH_1; // @[Bus.scala 265:25]
  wire  slaveMux_io_in_0_ready; // @[Bus.scala 310:26]
  wire  slaveMux_io_in_0_valid; // @[Bus.scala 310:26]
  wire [2:0] slaveMux_io_in_0_bits_opcode; // @[Bus.scala 310:26]
  wire [127:0] slaveMux_io_in_0_bits_data; // @[Bus.scala 310:26]
  wire  slaveMux_io_out_ready; // @[Bus.scala 310:26]
  wire  slaveMux_io_out_valid; // @[Bus.scala 310:26]
  wire [2:0] slaveMux_io_out_bits_opcode; // @[Bus.scala 310:26]
  wire [127:0] slaveMux_io_out_bits_data; // @[Bus.scala 310:26]
  wire  slaveMux_io_choseOH_0; // @[Bus.scala 310:26]
  wire [1:0] _WIRE_1 = reqArb_io_grantOH; // @[Bus.scala 238:{52,52}]
  reg  s1_full; // @[Bus.scala 249:26]
  wire  s1_latch = buf__io_deq_ready & buf__io_deq_valid; // @[Decoupled.scala 51:35]
  reg [2:0] s1_req_opcode; // @[Reg.scala 19:16]
  reg [127:0] s1_req_size; // @[Reg.scala 19:16]
  reg  s1_req_source; // @[Reg.scala 19:16]
  reg [31:0] s1_req_address; // @[Reg.scala 19:16]
  reg [127:0] s1_req_data; // @[Reg.scala 19:16]
  wire [123:0] s1_beatSize = s1_req_size[127:4]; // @[Bus.scala 255:35]
  reg [4:0] s1_beatCounter_value; // @[Counter.scala 61:40]
  wire [123:0] _s1_lastBeat_T_1 = s1_beatSize - 124'h1; // @[Bus.scala 278:60]
  wire [123:0] _GEN_27 = {{119'd0}, s1_beatCounter_value}; // @[Bus.scala 278:44]
  wire  s1_lastBeat = _GEN_27 == _s1_lastBeat_T_1; // @[Bus.scala 278:44]
  wire  _s1_putMultiBeat_T = ~s1_lastBeat; // @[Bus.scala 287:25]
  wire  _s1_putMultiBeat_T_1 = s1_req_opcode == 3'h2; // @[Bus.scala 287:55]
  wire  s1_putMultiBeat = ~s1_lastBeat & s1_req_opcode == 3'h2; // @[Bus.scala 287:38]
  reg  s2_full; // @[Bus.scala 297:26]
  reg [2:0] s2_opcode; // @[Reg.scala 19:16]
  wire [1:0] s2_masterRecvVec = {io_masterFace_out_1_valid,io_masterFace_out_0_valid}; // @[Cat.scala 33:92]
  reg [1:0] s2_chosenMasterOH; // @[Reg.scala 19:16]
  wire [1:0] _s2_masterRecv_T = s2_masterRecvVec & s2_chosenMasterOH; // @[Bus.scala 322:43]
  wire  s2_masterRecv = |_s2_masterRecv_T; // @[Bus.scala 322:64]
  reg  s2_masterRecvHold_holdReg; // @[Reg.scala 19:16]
  wire  s2_masterRecvHold = s2_masterRecv ? s2_masterRecv : s2_masterRecvHold_holdReg; // @[util.scala 26:12]
  reg [4:0] s2_beatCounter_value; // @[Counter.scala 61:40]
  reg [123:0] s2_beatSize; // @[Reg.scala 19:16]
  wire [123:0] _s2_lastBeat_T_1 = s2_beatSize - 124'h1; // @[Bus.scala 324:60]
  wire [123:0] _GEN_28 = {{119'd0}, s2_beatCounter_value}; // @[Bus.scala 324:44]
  wire  s2_lastBeat = _GEN_28 == _s2_lastBeat_T_1; // @[Bus.scala 324:44]
  wire  s2_getAllBeat = s2_opcode == 3'h4 & s2_masterRecvHold & s2_lastBeat; // @[Bus.scala 332:61]
  wire  s2_fire = s2_opcode == 3'h2 & s2_masterRecvHold | s2_getAllBeat; // @[Bus.scala 333:65]
  wire  s2_ready = ~s2_full | s2_fire; // @[Bus.scala 306:26]
  wire  _s1_slaveRecVec_T = io_slaveFace_in_0_ready & io_slaveFace_in_0_valid; // @[Decoupled.scala 51:35]
  wire [1:0] s1_slaveRecVec = {1'h0,_s1_slaveRecVec_T}; // @[Cat.scala 33:92]
  wire [1:0] _s1_slaveRecv_T = {addrDec_io_choseOH_1,addrDec_io_choseOH_0}; // @[Bus.scala 276:59]
  wire [1:0] _s1_slaveRecv_T_1 = s1_slaveRecVec & _s1_slaveRecv_T; // @[Bus.scala 276:40]
  wire  s1_slaveRecv = |_s1_slaveRecv_T_1; // @[Bus.scala 276:67]
  reg  s1_slaveRecvHold_holdReg; // @[Reg.scala 19:16]
  wire  s1_slaveRecvHold = s1_slaveRecv ? s1_slaveRecv : s1_slaveRecvHold_holdReg; // @[util.scala 26:12]
  wire  s1_putAllBeat = s1_lastBeat & _s1_putMultiBeat_T_1; // @[Bus.scala 289:34]
  wire  s1_valid = s1_slaveRecvHold & (s1_putAllBeat | s1_req_opcode == 3'h4); // @[Bus.scala 290:34]
  wire  s1_fire = s2_ready & s1_valid; // @[Bus.scala 292:25]
  wire  _GEN_8 = s1_full & s1_fire ? 1'h0 : s1_full; // @[Bus.scala 249:26 263:{35,45}]
  wire  _GEN_9 = s1_latch | _GEN_8; // @[Bus.scala 262:{20,30}]
  wire [4:0] _value_T_1 = s1_beatCounter_value + 5'h1; // @[Counter.scala 77:24]
  reg  s2_chosenSlaveOH_0; // @[Reg.scala 19:16]
  wire [1:0] _s2_chosenMasterOH_T = 2'h1 << s1_req_source; // @[OneHot.scala 57:35]
  wire  _GEN_19 = s2_full & s2_fire ? 1'h0 : s2_full; // @[Bus.scala 297:26 308:{35,45}]
  wire  _GEN_20 = s1_fire | _GEN_19; // @[Bus.scala 307:{20,30}]
  wire [4:0] _value_T_3 = s2_beatCounter_value + 5'h1; // @[Counter.scala 77:24]
  reg  idle; // @[Bus.scala 337:23]
  wire  _GEN_25 = s2_fire | idle; // @[Bus.scala 341:26 342:14 337:23]
  wire  _GEN_26 = s1_latch | s1_fire ? 1'h0 : _GEN_25; // @[Bus.scala 339:32 340:14]
  TLBusArbiter reqArb ( // @[Bus.scala 233:24]
    .clock(reqArb_clock),
    .reset(reqArb_reset),
    .io_reqs_1(reqArb_io_reqs_1),
    .io_grantOH(reqArb_io_grantOH)
  );
  TLBusMux reqMux ( // @[Bus.scala 236:24]
    .io_in_0_ready(reqMux_io_in_0_ready),
    .io_in_0_valid(reqMux_io_in_0_valid),
    .io_in_0_bits_address(reqMux_io_in_0_bits_address),
    .io_in_1_ready(reqMux_io_in_1_ready),
    .io_in_1_valid(reqMux_io_in_1_valid),
    .io_in_1_bits_opcode(reqMux_io_in_1_bits_opcode),
    .io_in_1_bits_address(reqMux_io_in_1_bits_address),
    .io_in_1_bits_data(reqMux_io_in_1_bits_data),
    .io_out_ready(reqMux_io_out_ready),
    .io_out_valid(reqMux_io_out_valid),
    .io_out_bits_opcode(reqMux_io_out_bits_opcode),
    .io_out_bits_size(reqMux_io_out_bits_size),
    .io_out_bits_source(reqMux_io_out_bits_source),
    .io_out_bits_address(reqMux_io_out_bits_address),
    .io_out_bits_data(reqMux_io_out_bits_data),
    .io_choseOH_0(reqMux_io_choseOH_0),
    .io_choseOH_1(reqMux_io_choseOH_1)
  );
  Queue_6 buf_ ( // @[Bus.scala 242:21]
    .clock(buf__clock),
    .reset(buf__reset),
    .io_enq_ready(buf__io_enq_ready),
    .io_enq_valid(buf__io_enq_valid),
    .io_enq_bits_opcode(buf__io_enq_bits_opcode),
    .io_enq_bits_size(buf__io_enq_bits_size),
    .io_enq_bits_source(buf__io_enq_bits_source),
    .io_enq_bits_address(buf__io_enq_bits_address),
    .io_enq_bits_data(buf__io_enq_bits_data),
    .io_deq_ready(buf__io_deq_ready),
    .io_deq_valid(buf__io_deq_valid),
    .io_deq_bits_opcode(buf__io_deq_bits_opcode),
    .io_deq_bits_size(buf__io_deq_bits_size),
    .io_deq_bits_source(buf__io_deq_bits_source),
    .io_deq_bits_address(buf__io_deq_bits_address),
    .io_deq_bits_data(buf__io_deq_bits_data)
  );
  TLAddrDecode addrDec ( // @[Bus.scala 265:25]
    .io_addr(addrDec_io_addr),
    .io_choseOH_0(addrDec_io_choseOH_0),
    .io_choseOH_1(addrDec_io_choseOH_1)
  );
  TLBusMux_1 slaveMux ( // @[Bus.scala 310:26]
    .io_in_0_ready(slaveMux_io_in_0_ready),
    .io_in_0_valid(slaveMux_io_in_0_valid),
    .io_in_0_bits_opcode(slaveMux_io_in_0_bits_opcode),
    .io_in_0_bits_data(slaveMux_io_in_0_bits_data),
    .io_out_ready(slaveMux_io_out_ready),
    .io_out_valid(slaveMux_io_out_valid),
    .io_out_bits_opcode(slaveMux_io_out_bits_opcode),
    .io_out_bits_data(slaveMux_io_out_bits_data),
    .io_choseOH_0(slaveMux_io_choseOH_0)
  );
  assign io_masterFace_in_0_ready = reqMux_io_in_0_ready; // @[Bus.scala 237:58]
  assign io_masterFace_in_1_ready = reqMux_io_in_1_ready; // @[Bus.scala 237:58]
  assign io_masterFace_out_0_valid = slaveMux_io_out_valid & s2_chosenMasterOH[0]; // @[Bus.scala 316:43]
  assign io_masterFace_out_0_bits_opcode = slaveMux_io_out_bits_opcode; // @[Bus.scala 315:17]
  assign io_masterFace_out_0_bits_data = slaveMux_io_out_bits_data; // @[Bus.scala 315:17]
  assign io_masterFace_out_1_valid = slaveMux_io_out_valid & s2_chosenMasterOH[1]; // @[Bus.scala 316:43]
  assign io_masterFace_out_1_bits_opcode = slaveMux_io_out_bits_opcode; // @[Bus.scala 315:17]
  assign io_masterFace_out_1_bits_data = slaveMux_io_out_bits_data; // @[Bus.scala 315:17]
  assign io_slaveFace_in_0_valid = addrDec_io_choseOH_0 & s1_full; // @[Bus.scala 271:41]
  assign io_slaveFace_in_0_bits_opcode = s1_req_opcode; // @[Bus.scala 270:18]
  assign io_slaveFace_in_0_bits_size = s1_req_size; // @[Bus.scala 270:18]
  assign io_slaveFace_in_0_bits_address = s1_req_address; // @[Bus.scala 270:18]
  assign io_slaveFace_in_0_bits_data = s1_req_data; // @[Bus.scala 270:18]
  assign io_slaveFace_out_0_ready = slaveMux_io_in_0_ready; // @[Bus.scala 311:20]
  assign reqArb_clock = clock;
  assign reqArb_reset = reset;
  assign reqArb_io_reqs_1 = io_masterFace_in_1_valid; // @[Bus.scala 234:58]
  assign reqMux_io_in_0_valid = io_masterFace_in_0_valid; // @[Bus.scala 237:58]
  assign reqMux_io_in_0_bits_address = io_masterFace_in_0_bits_address; // @[Bus.scala 237:58]
  assign reqMux_io_in_1_valid = io_masterFace_in_1_valid; // @[Bus.scala 237:58]
  assign reqMux_io_in_1_bits_opcode = io_masterFace_in_1_bits_opcode; // @[Bus.scala 237:58]
  assign reqMux_io_in_1_bits_address = io_masterFace_in_1_bits_address; // @[Bus.scala 237:58]
  assign reqMux_io_in_1_bits_data = io_masterFace_in_1_bits_data; // @[Bus.scala 237:58]
  assign reqMux_io_out_ready = buf__io_enq_ready; // @[Bus.scala 243:16]
  assign reqMux_io_choseOH_0 = _WIRE_1[0]; // @[Bus.scala 238:52]
  assign reqMux_io_choseOH_1 = _WIRE_1[1]; // @[Bus.scala 238:52]
  assign buf__clock = clock;
  assign buf__reset = reset;
  assign buf__io_enq_valid = reqMux_io_out_valid; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_opcode = reqMux_io_out_bits_opcode; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_size = reqMux_io_out_bits_size; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_source = reqMux_io_out_bits_source; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_address = reqMux_io_out_bits_address; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_data = reqMux_io_out_bits_data; // @[Bus.scala 243:16]
  assign buf__io_deq_ready = ~s1_full | s1_putMultiBeat | s1_fire; // @[Bus.scala 261:45]
  assign addrDec_io_addr = s1_req_address; // @[Bus.scala 267:21]
  assign slaveMux_io_in_0_valid = io_slaveFace_out_0_valid; // @[Bus.scala 311:20]
  assign slaveMux_io_in_0_bits_opcode = io_slaveFace_out_0_bits_opcode; // @[Bus.scala 311:20]
  assign slaveMux_io_in_0_bits_data = io_slaveFace_out_0_bits_data; // @[Bus.scala 311:20]
  assign slaveMux_io_out_ready = s2_chosenMasterOH[0] | s2_chosenMasterOH[1]; // @[Mux.scala 27:73]
  assign slaveMux_io_choseOH_0 = s2_chosenSlaveOH_0; // @[Bus.scala 312:25]
  always @(posedge clock) begin
    if (reset) begin // @[Bus.scala 249:26]
      s1_full <= 1'h0; // @[Bus.scala 249:26]
    end else begin
      s1_full <= _GEN_9;
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_opcode <= buf__io_deq_bits_opcode; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_size <= buf__io_deq_bits_size; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_source <= buf__io_deq_bits_source; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_address <= buf__io_deq_bits_address; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_data <= buf__io_deq_bits_data; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Counter.scala 61:40]
      s1_beatCounter_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (s1_fire) begin // @[Bus.scala 282:19]
      s1_beatCounter_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (s1_slaveRecv & _s1_putMultiBeat_T) begin // @[Bus.scala 279:40]
      s1_beatCounter_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Bus.scala 297:26]
      s2_full <= 1'h0; // @[Bus.scala 297:26]
    end else begin
      s2_full <= _GEN_20;
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_opcode <= s1_req_opcode; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_chosenMasterOH <= _s2_chosenMasterOH_T; // @[Reg.scala 20:22]
    end
    if (s2_fire) begin // @[util.scala 25:21]
      s2_masterRecvHold_holdReg <= 1'h0; // @[util.scala 25:31]
    end else if (s2_masterRecv) begin // @[util.scala 26:12]
      s2_masterRecvHold_holdReg <= s2_masterRecv;
    end
    if (reset) begin // @[Counter.scala 61:40]
      s2_beatCounter_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (s2_fire) begin // @[Bus.scala 328:19]
      s2_beatCounter_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (s2_masterRecv & ~s2_lastBeat) begin // @[Bus.scala 325:41]
      s2_beatCounter_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_beatSize <= s1_beatSize; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[util.scala 25:21]
      s1_slaveRecvHold_holdReg <= 1'h0; // @[util.scala 25:31]
    end else if (s1_slaveRecv) begin // @[util.scala 26:12]
      s1_slaveRecvHold_holdReg <= s1_slaveRecv;
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_chosenSlaveOH_0 <= addrDec_io_choseOH_0; // @[Reg.scala 20:22]
    end
    idle <= reset | _GEN_26; // @[Bus.scala 337:{23,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s1_req_opcode = _RAND_1[2:0];
  _RAND_2 = {4{`RANDOM}};
  s1_req_size = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  s1_req_source = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s1_req_address = _RAND_4[31:0];
  _RAND_5 = {4{`RANDOM}};
  s1_req_data = _RAND_5[127:0];
  _RAND_6 = {1{`RANDOM}};
  s1_beatCounter_value = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  s2_full = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s2_opcode = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  s2_chosenMasterOH = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  s2_masterRecvHold_holdReg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  s2_beatCounter_value = _RAND_11[4:0];
  _RAND_12 = {4{`RANDOM}};
  s2_beatSize = _RAND_12[123:0];
  _RAND_13 = {1{`RANDOM}};
  s1_slaveRecvHold_holdReg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  s2_chosenSlaveOH_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  idle = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SingleROM(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [2:0]   io_req_bits_opcode,
  input  [127:0] io_req_bits_size,
  input  [31:0]  io_req_bits_address,
  input  [127:0] io_req_bits_data,
  input          io_resp_ready,
  output         io_resp_valid,
  output [2:0]   io_resp_bits_opcode,
  output [127:0] io_resp_bits_size,
  output [127:0] io_resp_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] mem [0:131071]; // @[SingleROM.scala 14:26]
  wire  mem_rdata_en; // @[SingleROM.scala 14:26]
  wire [16:0] mem_rdata_addr; // @[SingleROM.scala 14:26]
  wire [127:0] mem_rdata_data; // @[SingleROM.scala 14:26]
  wire [127:0] mem_MPORT_data; // @[SingleROM.scala 14:26]
  wire [16:0] mem_MPORT_addr; // @[SingleROM.scala 14:26]
  wire  mem_MPORT_mask; // @[SingleROM.scala 14:26]
  wire  mem_MPORT_en; // @[SingleROM.scala 14:26]
  reg  mem_rdata_en_pipe_0;
  reg [16:0] mem_rdata_addr_pipe_0;
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [2:0] reqReg_opcode; // @[Reg.scala 19:16]
  reg [127:0] reqReg_size; // @[Reg.scala 19:16]
  reg [31:0] reqReg_address; // @[Reg.scala 19:16]
  reg [127:0] reqReg_data; // @[Reg.scala 19:16]
  wire [2:0] _GEN_0 = _reqReg_T ? io_req_bits_opcode : reqReg_opcode; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_4 = _reqReg_T ? io_req_bits_address : reqReg_address; // @[Reg.scala 19:16 20:{18,22}]
  reg  busy; // @[SingleROM.scala 19:23]
  reg [4:0] reqLastBeat_count_value; // @[Counter.scala 61:40]
  wire [123:0] reqLastBeat_beatNum = io_req_bits_size[127:4]; // @[Bus.scala 85:41]
  wire [123:0] _reqLastBeat_lastBeat_T_1 = reqLastBeat_beatNum - 124'h1; // @[Bus.scala 86:52]
  wire [123:0] _GEN_25 = {{119'd0}, reqLastBeat_count_value}; // @[Bus.scala 86:40]
  wire  reqLastBeat_lastBeat = _GEN_25 == _reqLastBeat_lastBeat_T_1; // @[Bus.scala 86:40]
  wire  reqLastBeat_fireLastBeat = _reqReg_T & reqLastBeat_lastBeat; // @[Bus.scala 87:38]
  wire [4:0] _reqLastBeat_value_T_1 = reqLastBeat_count_value + 5'h1; // @[Counter.scala 77:24]
  reg [4:0] respLastBeat_count_value; // @[Counter.scala 61:40]
  wire [123:0] respLastBeat_beatNum = io_resp_bits_size[127:4]; // @[Bus.scala 96:42]
  wire [123:0] _respLastBeat_lastBeat_T_1 = respLastBeat_beatNum - 124'h1; // @[Bus.scala 97:52]
  wire [123:0] _GEN_26 = {{119'd0}, respLastBeat_count_value}; // @[Bus.scala 97:40]
  wire  respLastBeat_lastBeat = _GEN_26 == _respLastBeat_lastBeat_T_1; // @[Bus.scala 97:40]
  wire  _respLastBeat_fireLastBeat_T = io_resp_ready & io_resp_valid; // @[Decoupled.scala 51:35]
  wire  respLastBeat_fireLastBeat = _respLastBeat_fireLastBeat_T & respLastBeat_lastBeat; // @[Bus.scala 98:39]
  wire [4:0] _respLastBeat_value_T_1 = respLastBeat_count_value + 5'h1; // @[Counter.scala 77:24]
  wire  _getFire_T_1 = _GEN_0 == 3'h4; // @[SingleROM.scala 27:45]
  wire  getFire = _reqReg_T & _GEN_0 == 3'h4; // @[SingleROM.scala 27:31]
  wire  _putFire_T_2 = _GEN_0 == 3'h2; // @[SingleROM.scala 28:60]
  wire  putFire = _reqReg_T & reqLastBeat_fireLastBeat & _GEN_0 == 3'h2; // @[SingleROM.scala 28:46]
  wire  reqLatch = getFire | putFire; // @[SingleROM.scala 29:28]
  wire  _finish_T_2 = reqReg_opcode == 3'h4; // @[SingleROM.scala 58:86]
  wire  finish = _respLastBeat_fireLastBeat_T & (reqReg_opcode == 3'h2 | reqReg_opcode == 3'h4 &
    respLastBeat_fireLastBeat); // @[SingleROM.scala 58:28]
  wire  _GEN_12 = busy & finish ? 1'h0 : busy; // @[SingleROM.scala 19:23 31:{31,38}]
  wire  _GEN_13 = reqLatch | _GEN_12; // @[SingleROM.scala 30:{20,27}]
  wire  ren = _getFire_T_1 & (_reqReg_T | _respLastBeat_fireLastBeat_T); // @[SingleROM.scala 33:41]
  wire  wen = _reqReg_T & _putFire_T_2; // @[SingleROM.scala 34:27]
  reg [4:0] beatCount_count_value; // @[Counter.scala 61:40]
  wire [123:0] _GEN_27 = {{119'd0}, beatCount_count_value}; // @[Bus.scala 97:40]
  wire  beatCount_lastBeat = _GEN_27 == _respLastBeat_lastBeat_T_1; // @[Bus.scala 97:40]
  wire  beatCount_fireLastBeat = _respLastBeat_fireLastBeat_T & beatCount_lastBeat; // @[Bus.scala 98:39]
  wire [4:0] _beatCount_value_T_1 = beatCount_count_value + 5'h1; // @[Counter.scala 77:24]
  wire [4:0] beatCount = _reqReg_T ? 5'h0 : _beatCount_value_T_1; // @[SingleROM.scala 38:24]
  wire [8:0] addrOff = {beatCount, 4'h0}; // @[SingleROM.scala 39:29]
  wire [31:0] _GEN_28 = {{23'd0}, addrOff}; // @[SingleROM.scala 40:31]
  wire [31:0] _rdAddr_T_1 = _GEN_4 + _GEN_28; // @[SingleROM.scala 40:31]
  wire [27:0] rdAddr = _rdAddr_T_1[31:4]; // @[SingleROM.scala 40:42]
  wire [27:0] wrAddr = _GEN_4[31:4]; // @[SingleROM.scala 45:30]
  assign mem_rdata_en = mem_rdata_en_pipe_0;
  assign mem_rdata_addr = mem_rdata_addr_pipe_0;
  assign mem_rdata_data = mem[mem_rdata_addr]; // @[SingleROM.scala 14:26]
  assign mem_MPORT_data = _reqReg_T ? io_req_bits_data : reqReg_data;
  assign mem_MPORT_addr = wrAddr[16:0];
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = wen;
  assign io_req_ready = ~busy; // @[SingleROM.scala 22:21]
  assign io_resp_valid = busy; // @[SingleROM.scala 51:19]
  assign io_resp_bits_opcode = {{2'd0}, _finish_T_2}; // @[SingleROM.scala 55:25]
  assign io_resp_bits_size = reqReg_size; // @[SingleROM.scala 53:23]
  assign io_resp_bits_data = mem_rdata_data; // @[SingleROM.scala 54:23]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SingleROM.scala 14:26]
    end
    mem_rdata_en_pipe_0 <= ren;
    if (ren) begin
      mem_rdata_addr_pipe_0 <= rdAddr[16:0];
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_opcode <= io_req_bits_opcode; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_size <= io_req_bits_size; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_address <= io_req_bits_address; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data <= io_req_bits_data; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[SingleROM.scala 19:23]
      busy <= 1'h0; // @[SingleROM.scala 19:23]
    end else begin
      busy <= _GEN_13;
    end
    if (reset) begin // @[Counter.scala 61:40]
      reqLastBeat_count_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (reqLastBeat_fireLastBeat | _reqReg_T & io_req_bits_opcode == 3'h4) begin // @[Bus.scala 88:71]
      reqLastBeat_count_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (_reqReg_T) begin // @[Bus.scala 90:34]
      reqLastBeat_count_value <= _reqLastBeat_value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      respLastBeat_count_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (respLastBeat_fireLastBeat | _respLastBeat_fireLastBeat_T & io_resp_bits_opcode == 3'h0) begin // @[Bus.scala 99:79]
      respLastBeat_count_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (_respLastBeat_fireLastBeat_T) begin // @[Bus.scala 101:35]
      respLastBeat_count_value <= _respLastBeat_value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      beatCount_count_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (beatCount_fireLastBeat | _respLastBeat_fireLastBeat_T & io_resp_bits_opcode == 3'h0) begin // @[Bus.scala 99:79]
      beatCount_count_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (_respLastBeat_fireLastBeat_T) begin // @[Bus.scala 101:35]
      beatCount_count_value <= _beatCount_value_T_1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 131072; initvar = initvar+1)
    mem[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_rdata_addr_pipe_0 = _RAND_2[16:0];
  _RAND_3 = {1{`RANDOM}};
  reqReg_opcode = _RAND_3[2:0];
  _RAND_4 = {4{`RANDOM}};
  reqReg_size = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  reqReg_address = _RAND_5[31:0];
  _RAND_6 = {4{`RANDOM}};
  reqReg_data = _RAND_6[127:0];
  _RAND_7 = {1{`RANDOM}};
  busy = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reqLastBeat_count_value = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  respLastBeat_count_value = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  beatCount_count_value = _RAND_10[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  input         io_in_start,
  output [31:0] io_out_state_intRegState_regState_0,
  output [31:0] io_out_state_intRegState_regState_1,
  output [31:0] io_out_state_intRegState_regState_2,
  output [31:0] io_out_state_intRegState_regState_3,
  output [31:0] io_out_state_intRegState_regState_4,
  output [31:0] io_out_state_intRegState_regState_5,
  output [31:0] io_out_state_intRegState_regState_6,
  output [31:0] io_out_state_intRegState_regState_7,
  output [31:0] io_out_state_intRegState_regState_8,
  output [31:0] io_out_state_intRegState_regState_9,
  output [31:0] io_out_state_intRegState_regState_10,
  output [31:0] io_out_state_intRegState_regState_11,
  output [31:0] io_out_state_intRegState_regState_12,
  output [31:0] io_out_state_intRegState_regState_13,
  output [31:0] io_out_state_intRegState_regState_14,
  output [31:0] io_out_state_intRegState_regState_15,
  output [31:0] io_out_state_intRegState_regState_16,
  output [31:0] io_out_state_intRegState_regState_17,
  output [31:0] io_out_state_intRegState_regState_18,
  output [31:0] io_out_state_intRegState_regState_19,
  output [31:0] io_out_state_intRegState_regState_20,
  output [31:0] io_out_state_intRegState_regState_21,
  output [31:0] io_out_state_intRegState_regState_22,
  output [31:0] io_out_state_intRegState_regState_23,
  output [31:0] io_out_state_intRegState_regState_24,
  output [31:0] io_out_state_intRegState_regState_25,
  output [31:0] io_out_state_intRegState_regState_26,
  output [31:0] io_out_state_intRegState_regState_27,
  output [31:0] io_out_state_intRegState_regState_28,
  output [31:0] io_out_state_intRegState_regState_29,
  output [31:0] io_out_state_intRegState_regState_30,
  output [31:0] io_out_state_intRegState_regState_31,
  output        io_out_state_instState_commit,
  output [31:0] io_out_state_instState_pc,
  output [31:0] io_out_state_instState_inst,
  output [31:0] io_out_state_csrState_mcycle,
  output [31:0] io_out_state_csrState_mcycleh
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
`endif // RANDOMIZE_REG_INIT
  wire  ib_clock; // @[Core_1.scala 50:20]
  wire  ib_reset; // @[Core_1.scala 50:20]
  wire  ib_io_in_ready; // @[Core_1.scala 50:20]
  wire  ib_io_in_valid; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_in_bits_icache_data; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_in_bits_icache_addr; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_in_bits_icache_inst_0; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_in_bits_icache_inst_1; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_in_bits_icache_inst_2; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_in_bits_icache_inst_3; // @[Core_1.scala 50:20]
  wire [2:0] ib_io_in_bits_icache_size; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_in_bits_pc; // @[Core_1.scala 50:20]
  wire  ib_io_in_bits_flush; // @[Core_1.scala 50:20]
  wire  ib_io_out_ready; // @[Core_1.scala 50:20]
  wire  ib_io_out_valid; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_out_bits_inst_0_inst; // @[Core_1.scala 50:20]
  wire  ib_io_out_bits_inst_0_valid; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_out_bits_inst_1_inst; // @[Core_1.scala 50:20]
  wire  ib_io_out_bits_inst_1_valid; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_out_bits_inst_2_inst; // @[Core_1.scala 50:20]
  wire  ib_io_out_bits_inst_2_valid; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_out_bits_inst_3_inst; // @[Core_1.scala 50:20]
  wire  ib_io_out_bits_inst_3_valid; // @[Core_1.scala 50:20]
  wire [31:0] ib_io_out_bits_pc; // @[Core_1.scala 50:20]
  wire  ib_io_status_back_pressure; // @[Core_1.scala 50:20]
  wire  ib_io_status_full; // @[Core_1.scala 50:20]
  wire  icache_clock; // @[Core_1.scala 52:24]
  wire  icache_reset; // @[Core_1.scala 52:24]
  wire  icache_io_read_req_ready; // @[Core_1.scala 52:24]
  wire  icache_io_read_req_valid; // @[Core_1.scala 52:24]
  wire [31:0] icache_io_read_req_bits_addr; // @[Core_1.scala 52:24]
  wire  icache_io_read_resp_ready; // @[Core_1.scala 52:24]
  wire  icache_io_read_resp_valid; // @[Core_1.scala 52:24]
  wire [31:0] icache_io_read_resp_bits_data; // @[Core_1.scala 52:24]
  wire [31:0] icache_io_read_resp_bits_addr; // @[Core_1.scala 52:24]
  wire [31:0] icache_io_read_resp_bits_inst_0; // @[Core_1.scala 52:24]
  wire [31:0] icache_io_read_resp_bits_inst_1; // @[Core_1.scala 52:24]
  wire [31:0] icache_io_read_resp_bits_inst_2; // @[Core_1.scala 52:24]
  wire [31:0] icache_io_read_resp_bits_inst_3; // @[Core_1.scala 52:24]
  wire [2:0] icache_io_read_resp_bits_size; // @[Core_1.scala 52:24]
  wire  icache_io_tlbus_req_ready; // @[Core_1.scala 52:24]
  wire  icache_io_tlbus_req_valid; // @[Core_1.scala 52:24]
  wire [31:0] icache_io_tlbus_req_bits_address; // @[Core_1.scala 52:24]
  wire  icache_io_tlbus_resp_ready; // @[Core_1.scala 52:24]
  wire  icache_io_tlbus_resp_valid; // @[Core_1.scala 52:24]
  wire [2:0] icache_io_tlbus_resp_bits_opcode; // @[Core_1.scala 52:24]
  wire [127:0] icache_io_tlbus_resp_bits_data; // @[Core_1.scala 52:24]
  wire  icache_io_flush; // @[Core_1.scala 52:24]
  wire  rf_clock; // @[Core_1.scala 64:20]
  wire  rf_reset; // @[Core_1.scala 64:20]
  wire [4:0] rf_io_r_0_addr; // @[Core_1.scala 64:20]
  wire [31:0] rf_io_r_0_data; // @[Core_1.scala 64:20]
  wire [4:0] rf_io_r_1_addr; // @[Core_1.scala 64:20]
  wire [31:0] rf_io_r_1_data; // @[Core_1.scala 64:20]
  wire [4:0] rf_io_r_2_addr; // @[Core_1.scala 64:20]
  wire [31:0] rf_io_r_2_data; // @[Core_1.scala 64:20]
  wire [4:0] rf_io_r_3_addr; // @[Core_1.scala 64:20]
  wire [31:0] rf_io_r_3_data; // @[Core_1.scala 64:20]
  wire [4:0] rf_io_r_4_addr; // @[Core_1.scala 64:20]
  wire [31:0] rf_io_r_4_data; // @[Core_1.scala 64:20]
  wire [4:0] rf_io_r_5_addr; // @[Core_1.scala 64:20]
  wire [31:0] rf_io_r_5_data; // @[Core_1.scala 64:20]
  wire [4:0] rf_io_r_6_addr; // @[Core_1.scala 64:20]
  wire [31:0] rf_io_r_6_data; // @[Core_1.scala 64:20]
  wire [4:0] rf_io_r_7_addr; // @[Core_1.scala 64:20]
  wire [31:0] rf_io_r_7_data; // @[Core_1.scala 64:20]
  wire [4:0] rf_io_w_0_addr; // @[Core_1.scala 64:20]
  wire  rf_io_w_0_en; // @[Core_1.scala 64:20]
  wire [31:0] rf_io_w_0_data; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_0; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_1; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_2; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_3; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_4; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_5; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_6; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_7; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_8; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_9; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_10; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_11; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_12; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_13; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_14; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_15; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_16; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_17; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_18; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_19; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_20; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_21; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_22; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_23; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_24; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_25; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_26; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_27; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_28; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_29; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_30; // @[Core_1.scala 64:20]
  wire [31:0] rf_regState_0_regState_31; // @[Core_1.scala 64:20]
  wire  rob_clock; // @[Core_1.scala 79:21]
  wire  rob_reset; // @[Core_1.scala 79:21]
  wire  rob_io_enq_ready; // @[Core_1.scala 79:21]
  wire  rob_io_enq_valid; // @[Core_1.scala 79:21]
  wire [4:0] rob_io_enq_bits_rd; // @[Core_1.scala 79:21]
  wire [3:0] rob_io_enq_bits_fuValid; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_enq_bits_fuOp; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_enq_bits_pc; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_enq_bits_inst; // @[Core_1.scala 79:21]
  wire  rob_io_deq_ready; // @[Core_1.scala 79:21]
  wire  rob_io_deq_valid; // @[Core_1.scala 79:21]
  wire  rob_io_deq_bits_rdWrEn; // @[Core_1.scala 79:21]
  wire [4:0] rob_io_deq_bits_rd; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_deq_bits_data; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_deq_bits_id; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_deq_bits_brAddr; // @[Core_1.scala 79:21]
  wire  rob_io_deq_bits_brTaken; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_deq_bits_excpAddr; // @[Core_1.scala 79:21]
  wire  rob_io_deq_bits_excpValid; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_deq_bits_pc; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_deq_bits_inst; // @[Core_1.scala 79:21]
  wire  rob_io_rs_0_valid; // @[Core_1.scala 79:21]
  wire [2:0] rob_io_rs_0_bits_id; // @[Core_1.scala 79:21]
  wire  rob_io_rs_1_valid; // @[Core_1.scala 79:21]
  wire [2:0] rob_io_rs_1_bits_id; // @[Core_1.scala 79:21]
  wire  rob_io_rs_2_valid; // @[Core_1.scala 79:21]
  wire [2:0] rob_io_rs_2_bits_id; // @[Core_1.scala 79:21]
  wire  rob_io_rs_3_valid; // @[Core_1.scala 79:21]
  wire [2:0] rob_io_rs_3_bits_id; // @[Core_1.scala 79:21]
  wire  rob_io_read_0_busy; // @[Core_1.scala 79:21]
  wire [1:0] rob_io_read_0_state; // @[Core_1.scala 79:21]
  wire [4:0] rob_io_read_0_rd; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_read_0_data; // @[Core_1.scala 79:21]
  wire  rob_io_read_1_busy; // @[Core_1.scala 79:21]
  wire [1:0] rob_io_read_1_state; // @[Core_1.scala 79:21]
  wire [4:0] rob_io_read_1_rd; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_read_1_data; // @[Core_1.scala 79:21]
  wire  rob_io_read_2_busy; // @[Core_1.scala 79:21]
  wire [1:0] rob_io_read_2_state; // @[Core_1.scala 79:21]
  wire [4:0] rob_io_read_2_rd; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_read_2_data; // @[Core_1.scala 79:21]
  wire  rob_io_read_3_busy; // @[Core_1.scala 79:21]
  wire [1:0] rob_io_read_3_state; // @[Core_1.scala 79:21]
  wire [4:0] rob_io_read_3_rd; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_read_3_data; // @[Core_1.scala 79:21]
  wire  rob_io_read_4_busy; // @[Core_1.scala 79:21]
  wire [1:0] rob_io_read_4_state; // @[Core_1.scala 79:21]
  wire [4:0] rob_io_read_4_rd; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_read_4_data; // @[Core_1.scala 79:21]
  wire  rob_io_fu_0_valid; // @[Core_1.scala 79:21]
  wire [2:0] rob_io_fu_0_bits_id; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_fu_0_bits_data; // @[Core_1.scala 79:21]
  wire  rob_io_fu_1_valid; // @[Core_1.scala 79:21]
  wire [2:0] rob_io_fu_1_bits_id; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_fu_1_bits_data; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_fu_1_bits_brAddr; // @[Core_1.scala 79:21]
  wire  rob_io_fu_1_bits_brTaken; // @[Core_1.scala 79:21]
  wire  rob_io_fu_2_valid; // @[Core_1.scala 79:21]
  wire [2:0] rob_io_fu_2_bits_id; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_fu_2_bits_data; // @[Core_1.scala 79:21]
  wire  rob_io_fu_3_valid; // @[Core_1.scala 79:21]
  wire [2:0] rob_io_fu_3_bits_id; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_fu_3_bits_data; // @[Core_1.scala 79:21]
  wire [31:0] rob_io_fu_3_bits_excpAddr; // @[Core_1.scala 79:21]
  wire  rob_io_fu_3_bits_excpValid; // @[Core_1.scala 79:21]
  wire [2:0] rob_io_id; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_0_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_1_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_2_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_3_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_4_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_5_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_6_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_7_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_8_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_9_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_10_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_11_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_12_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_13_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_14_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_15_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_16_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_17_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_18_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_19_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_20_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_21_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_22_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_23_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_24_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_25_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_26_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_27_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_28_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_29_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_30_owner; // @[Core_1.scala 79:21]
  wire [7:0] rob_io_regStatus_31_owner; // @[Core_1.scala 79:21]
  wire  rob_io_flush; // @[Core_1.scala 79:21]
  wire  aluStage_1_clock; // @[Core_1.scala 81:28]
  wire  aluStage_1_reset; // @[Core_1.scala 81:28]
  wire  aluStage_1_io_in_ready; // @[Core_1.scala 81:28]
  wire  aluStage_1_io_in_valid; // @[Core_1.scala 81:28]
  wire [3:0] aluStage_1_io_in_bits_opr1; // @[Core_1.scala 81:28]
  wire [3:0] aluStage_1_io_in_bits_opr2; // @[Core_1.scala 81:28]
  wire [4:0] aluStage_1_io_in_bits_aluOp; // @[Core_1.scala 81:28]
  wire [2:0] aluStage_1_io_in_bits_immSrc; // @[Core_1.scala 81:28]
  wire  aluStage_1_io_in_bits_immSign; // @[Core_1.scala 81:28]
  wire [31:0] aluStage_1_io_in_bits_rs1Val; // @[Core_1.scala 81:28]
  wire [31:0] aluStage_1_io_in_bits_rs2Val; // @[Core_1.scala 81:28]
  wire [31:0] aluStage_1_io_in_bits_inst; // @[Core_1.scala 81:28]
  wire [31:0] aluStage_1_io_in_bits_pc; // @[Core_1.scala 81:28]
  wire [7:0] aluStage_1_io_in_bits_id; // @[Core_1.scala 81:28]
  wire  aluStage_1_io_out_valid; // @[Core_1.scala 81:28]
  wire [31:0] aluStage_1_io_out_bits_data; // @[Core_1.scala 81:28]
  wire [7:0] aluStage_1_io_out_bits_id; // @[Core_1.scala 81:28]
  wire [4:0] aluStage_1_io_out_bits_rd; // @[Core_1.scala 81:28]
  wire  aluStage_1_io_flush; // @[Core_1.scala 81:28]
  wire  aluRS_clock; // @[Core_1.scala 82:23]
  wire  aluRS_reset; // @[Core_1.scala 82:23]
  wire  aluRS_io_enq_ready; // @[Core_1.scala 82:23]
  wire  aluRS_io_enq_valid; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_enq_bits_op; // @[Core_1.scala 82:23]
  wire [3:0] aluRS_io_enq_bits_opr1; // @[Core_1.scala 82:23]
  wire [3:0] aluRS_io_enq_bits_opr2; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_enq_bits_rs1; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_enq_bits_rs2; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_enq_bits_ROBId; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_enq_bits_rs1ROBId; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_enq_bits_rs2ROBId; // @[Core_1.scala 82:23]
  wire [2:0] aluRS_io_enq_bits_immSrc; // @[Core_1.scala 82:23]
  wire  aluRS_io_enq_bits_immSign; // @[Core_1.scala 82:23]
  wire [3:0] aluRS_io_enq_bits_excpType; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_enq_bits_pc; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_enq_bits_inst; // @[Core_1.scala 82:23]
  wire  aluRS_io_deq_ready; // @[Core_1.scala 82:23]
  wire  aluRS_io_deq_valid; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_deq_bits_op; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_deq_bits_ROBId; // @[Core_1.scala 82:23]
  wire [3:0] aluRS_io_deq_bits_opr1; // @[Core_1.scala 82:23]
  wire [3:0] aluRS_io_deq_bits_opr2; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_deq_bits_rs1Val; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_deq_bits_rs2Val; // @[Core_1.scala 82:23]
  wire [2:0] aluRS_io_deq_bits_immSrc; // @[Core_1.scala 82:23]
  wire  aluRS_io_deq_bits_immSign; // @[Core_1.scala 82:23]
  wire [3:0] aluRS_io_deq_bits_excpType; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_deq_bits_pc; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_deq_bits_inst; // @[Core_1.scala 82:23]
  wire  aluRS_io_robOut_valid; // @[Core_1.scala 82:23]
  wire [2:0] aluRS_io_robOut_bits_id; // @[Core_1.scala 82:23]
  wire  aluRS_io_robRead_0_busy; // @[Core_1.scala 82:23]
  wire [1:0] aluRS_io_robRead_0_state; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_robRead_0_rd; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_robRead_0_data; // @[Core_1.scala 82:23]
  wire  aluRS_io_robRead_1_busy; // @[Core_1.scala 82:23]
  wire [1:0] aluRS_io_robRead_1_state; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_robRead_1_rd; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_robRead_1_data; // @[Core_1.scala 82:23]
  wire  aluRS_io_robRead_2_busy; // @[Core_1.scala 82:23]
  wire [1:0] aluRS_io_robRead_2_state; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_robRead_2_rd; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_robRead_2_data; // @[Core_1.scala 82:23]
  wire  aluRS_io_robRead_3_busy; // @[Core_1.scala 82:23]
  wire [1:0] aluRS_io_robRead_3_state; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_robRead_3_rd; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_robRead_3_data; // @[Core_1.scala 82:23]
  wire  aluRS_io_robRead_4_busy; // @[Core_1.scala 82:23]
  wire [1:0] aluRS_io_robRead_4_state; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_robRead_4_rd; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_robRead_4_data; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_0_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_1_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_2_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_3_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_4_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_5_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_6_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_7_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_8_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_9_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_10_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_11_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_12_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_13_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_14_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_15_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_16_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_17_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_18_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_19_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_20_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_21_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_22_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_23_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_24_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_25_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_26_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_27_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_28_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_29_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_30_owner; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_regStatus_31_owner; // @[Core_1.scala 82:23]
  wire  aluRS_io_cdb_0_valid; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_cdb_0_bits_data; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_cdb_0_bits_id; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_cdb_0_bits_rd; // @[Core_1.scala 82:23]
  wire  aluRS_io_cdb_1_valid; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_cdb_1_bits_data; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_cdb_1_bits_id; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_cdb_1_bits_rd; // @[Core_1.scala 82:23]
  wire  aluRS_io_cdb_2_valid; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_cdb_2_bits_data; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_cdb_2_bits_id; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_cdb_2_bits_rd; // @[Core_1.scala 82:23]
  wire  aluRS_io_cdb_3_valid; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_cdb_3_bits_data; // @[Core_1.scala 82:23]
  wire [7:0] aluRS_io_cdb_3_bits_id; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_cdb_3_bits_rd; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_rf_0_addr; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_rf_0_data; // @[Core_1.scala 82:23]
  wire [4:0] aluRS_io_rf_1_addr; // @[Core_1.scala 82:23]
  wire [31:0] aluRS_io_rf_1_data; // @[Core_1.scala 82:23]
  wire  aluRS_io_flush; // @[Core_1.scala 82:23]
  wire  bruStage_1_clock; // @[Core_1.scala 84:28]
  wire  bruStage_1_reset; // @[Core_1.scala 84:28]
  wire  bruStage_1_io_in_ready; // @[Core_1.scala 84:28]
  wire  bruStage_1_io_in_valid; // @[Core_1.scala 84:28]
  wire [3:0] bruStage_1_io_in_bits_opr1; // @[Core_1.scala 84:28]
  wire [3:0] bruStage_1_io_in_bits_opr2; // @[Core_1.scala 84:28]
  wire [3:0] bruStage_1_io_in_bits_bruOp; // @[Core_1.scala 84:28]
  wire [2:0] bruStage_1_io_in_bits_immSrc; // @[Core_1.scala 84:28]
  wire [31:0] bruStage_1_io_in_bits_rs1Val; // @[Core_1.scala 84:28]
  wire [31:0] bruStage_1_io_in_bits_rs2Val; // @[Core_1.scala 84:28]
  wire [31:0] bruStage_1_io_in_bits_inst; // @[Core_1.scala 84:28]
  wire [31:0] bruStage_1_io_in_bits_pc; // @[Core_1.scala 84:28]
  wire [7:0] bruStage_1_io_in_bits_id; // @[Core_1.scala 84:28]
  wire  bruStage_1_io_out_valid; // @[Core_1.scala 84:28]
  wire  bruStage_1_io_out_bits_brTaken; // @[Core_1.scala 84:28]
  wire [31:0] bruStage_1_io_out_bits_brAddr; // @[Core_1.scala 84:28]
  wire [4:0] bruStage_1_io_out_bits_rd; // @[Core_1.scala 84:28]
  wire [31:0] bruStage_1_io_out_bits_data; // @[Core_1.scala 84:28]
  wire [7:0] bruStage_1_io_out_bits_id; // @[Core_1.scala 84:28]
  wire  bruStage_1_io_flush; // @[Core_1.scala 84:28]
  wire  bruRS_clock; // @[Core_1.scala 85:23]
  wire  bruRS_reset; // @[Core_1.scala 85:23]
  wire  bruRS_io_enq_ready; // @[Core_1.scala 85:23]
  wire  bruRS_io_enq_valid; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_enq_bits_op; // @[Core_1.scala 85:23]
  wire [3:0] bruRS_io_enq_bits_opr1; // @[Core_1.scala 85:23]
  wire [3:0] bruRS_io_enq_bits_opr2; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_enq_bits_rs1; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_enq_bits_rs2; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_enq_bits_ROBId; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_enq_bits_rs1ROBId; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_enq_bits_rs2ROBId; // @[Core_1.scala 85:23]
  wire [2:0] bruRS_io_enq_bits_immSrc; // @[Core_1.scala 85:23]
  wire  bruRS_io_enq_bits_immSign; // @[Core_1.scala 85:23]
  wire [3:0] bruRS_io_enq_bits_excpType; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_enq_bits_pc; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_enq_bits_inst; // @[Core_1.scala 85:23]
  wire  bruRS_io_deq_ready; // @[Core_1.scala 85:23]
  wire  bruRS_io_deq_valid; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_deq_bits_op; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_deq_bits_ROBId; // @[Core_1.scala 85:23]
  wire [3:0] bruRS_io_deq_bits_opr1; // @[Core_1.scala 85:23]
  wire [3:0] bruRS_io_deq_bits_opr2; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_deq_bits_rs1Val; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_deq_bits_rs2Val; // @[Core_1.scala 85:23]
  wire [2:0] bruRS_io_deq_bits_immSrc; // @[Core_1.scala 85:23]
  wire  bruRS_io_deq_bits_immSign; // @[Core_1.scala 85:23]
  wire [3:0] bruRS_io_deq_bits_excpType; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_deq_bits_pc; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_deq_bits_inst; // @[Core_1.scala 85:23]
  wire  bruRS_io_robOut_valid; // @[Core_1.scala 85:23]
  wire [2:0] bruRS_io_robOut_bits_id; // @[Core_1.scala 85:23]
  wire  bruRS_io_robRead_0_busy; // @[Core_1.scala 85:23]
  wire [1:0] bruRS_io_robRead_0_state; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_robRead_0_rd; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_robRead_0_data; // @[Core_1.scala 85:23]
  wire  bruRS_io_robRead_1_busy; // @[Core_1.scala 85:23]
  wire [1:0] bruRS_io_robRead_1_state; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_robRead_1_rd; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_robRead_1_data; // @[Core_1.scala 85:23]
  wire  bruRS_io_robRead_2_busy; // @[Core_1.scala 85:23]
  wire [1:0] bruRS_io_robRead_2_state; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_robRead_2_rd; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_robRead_2_data; // @[Core_1.scala 85:23]
  wire  bruRS_io_robRead_3_busy; // @[Core_1.scala 85:23]
  wire [1:0] bruRS_io_robRead_3_state; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_robRead_3_rd; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_robRead_3_data; // @[Core_1.scala 85:23]
  wire  bruRS_io_robRead_4_busy; // @[Core_1.scala 85:23]
  wire [1:0] bruRS_io_robRead_4_state; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_robRead_4_rd; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_robRead_4_data; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_0_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_1_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_2_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_3_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_4_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_5_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_6_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_7_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_8_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_9_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_10_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_11_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_12_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_13_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_14_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_15_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_16_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_17_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_18_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_19_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_20_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_21_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_22_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_23_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_24_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_25_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_26_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_27_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_28_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_29_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_30_owner; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_regStatus_31_owner; // @[Core_1.scala 85:23]
  wire  bruRS_io_cdb_0_valid; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_cdb_0_bits_data; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_cdb_0_bits_id; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_cdb_0_bits_rd; // @[Core_1.scala 85:23]
  wire  bruRS_io_cdb_1_valid; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_cdb_1_bits_data; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_cdb_1_bits_id; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_cdb_1_bits_rd; // @[Core_1.scala 85:23]
  wire  bruRS_io_cdb_2_valid; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_cdb_2_bits_data; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_cdb_2_bits_id; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_cdb_2_bits_rd; // @[Core_1.scala 85:23]
  wire  bruRS_io_cdb_3_valid; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_cdb_3_bits_data; // @[Core_1.scala 85:23]
  wire [7:0] bruRS_io_cdb_3_bits_id; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_cdb_3_bits_rd; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_rf_0_addr; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_rf_0_data; // @[Core_1.scala 85:23]
  wire [4:0] bruRS_io_rf_1_addr; // @[Core_1.scala 85:23]
  wire [31:0] bruRS_io_rf_1_data; // @[Core_1.scala 85:23]
  wire  bruRS_io_flush; // @[Core_1.scala 85:23]
  wire  lsuStage_1_clock; // @[Core_1.scala 87:28]
  wire  lsuStage_1_reset; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_in_ready; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_in_valid; // @[Core_1.scala 87:28]
  wire [4:0] lsuStage_1_io_in_bits_lsuOp; // @[Core_1.scala 87:28]
  wire [2:0] lsuStage_1_io_in_bits_immSrc; // @[Core_1.scala 87:28]
  wire [31:0] lsuStage_1_io_in_bits_rs1Val; // @[Core_1.scala 87:28]
  wire [31:0] lsuStage_1_io_in_bits_rs2Val; // @[Core_1.scala 87:28]
  wire [31:0] lsuStage_1_io_in_bits_inst; // @[Core_1.scala 87:28]
  wire [7:0] lsuStage_1_io_in_bits_id; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_out_valid; // @[Core_1.scala 87:28]
  wire [4:0] lsuStage_1_io_out_bits_rd; // @[Core_1.scala 87:28]
  wire [31:0] lsuStage_1_io_out_bits_data; // @[Core_1.scala 87:28]
  wire [7:0] lsuStage_1_io_out_bits_id; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_cache_read_req_ready; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_cache_read_req_valid; // @[Core_1.scala 87:28]
  wire [31:0] lsuStage_1_io_cache_read_req_bits_addr; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_cache_read_resp_ready; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_cache_read_resp_valid; // @[Core_1.scala 87:28]
  wire [31:0] lsuStage_1_io_cache_read_resp_bits_data; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_cache_write_req_ready; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_cache_write_req_valid; // @[Core_1.scala 87:28]
  wire [31:0] lsuStage_1_io_cache_write_req_bits_addr; // @[Core_1.scala 87:28]
  wire [31:0] lsuStage_1_io_cache_write_req_bits_data; // @[Core_1.scala 87:28]
  wire [3:0] lsuStage_1_io_cache_write_req_bits_mask; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_cache_write_resp_ready; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_cache_write_resp_valid; // @[Core_1.scala 87:28]
  wire [7:0] lsuStage_1_io_rob_bits_id; // @[Core_1.scala 87:28]
  wire  lsuStage_1_io_flush; // @[Core_1.scala 87:28]
  wire  lsuRS_clock; // @[Core_1.scala 88:23]
  wire  lsuRS_reset; // @[Core_1.scala 88:23]
  wire  lsuRS_io_enq_ready; // @[Core_1.scala 88:23]
  wire  lsuRS_io_enq_valid; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_enq_bits_op; // @[Core_1.scala 88:23]
  wire [3:0] lsuRS_io_enq_bits_opr1; // @[Core_1.scala 88:23]
  wire [3:0] lsuRS_io_enq_bits_opr2; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_enq_bits_rs1; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_enq_bits_rs2; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_enq_bits_ROBId; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_enq_bits_rs1ROBId; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_enq_bits_rs2ROBId; // @[Core_1.scala 88:23]
  wire [2:0] lsuRS_io_enq_bits_immSrc; // @[Core_1.scala 88:23]
  wire  lsuRS_io_enq_bits_immSign; // @[Core_1.scala 88:23]
  wire [3:0] lsuRS_io_enq_bits_excpType; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_enq_bits_pc; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_enq_bits_inst; // @[Core_1.scala 88:23]
  wire  lsuRS_io_deq_ready; // @[Core_1.scala 88:23]
  wire  lsuRS_io_deq_valid; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_deq_bits_op; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_deq_bits_ROBId; // @[Core_1.scala 88:23]
  wire [3:0] lsuRS_io_deq_bits_opr1; // @[Core_1.scala 88:23]
  wire [3:0] lsuRS_io_deq_bits_opr2; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_deq_bits_rs1Val; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_deq_bits_rs2Val; // @[Core_1.scala 88:23]
  wire [2:0] lsuRS_io_deq_bits_immSrc; // @[Core_1.scala 88:23]
  wire  lsuRS_io_deq_bits_immSign; // @[Core_1.scala 88:23]
  wire [3:0] lsuRS_io_deq_bits_excpType; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_deq_bits_pc; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_deq_bits_inst; // @[Core_1.scala 88:23]
  wire  lsuRS_io_robOut_valid; // @[Core_1.scala 88:23]
  wire [2:0] lsuRS_io_robOut_bits_id; // @[Core_1.scala 88:23]
  wire  lsuRS_io_robRead_0_busy; // @[Core_1.scala 88:23]
  wire [1:0] lsuRS_io_robRead_0_state; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_robRead_0_rd; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_robRead_0_data; // @[Core_1.scala 88:23]
  wire  lsuRS_io_robRead_1_busy; // @[Core_1.scala 88:23]
  wire [1:0] lsuRS_io_robRead_1_state; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_robRead_1_rd; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_robRead_1_data; // @[Core_1.scala 88:23]
  wire  lsuRS_io_robRead_2_busy; // @[Core_1.scala 88:23]
  wire [1:0] lsuRS_io_robRead_2_state; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_robRead_2_rd; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_robRead_2_data; // @[Core_1.scala 88:23]
  wire  lsuRS_io_robRead_3_busy; // @[Core_1.scala 88:23]
  wire [1:0] lsuRS_io_robRead_3_state; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_robRead_3_rd; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_robRead_3_data; // @[Core_1.scala 88:23]
  wire  lsuRS_io_robRead_4_busy; // @[Core_1.scala 88:23]
  wire [1:0] lsuRS_io_robRead_4_state; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_robRead_4_rd; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_robRead_4_data; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_0_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_1_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_2_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_3_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_4_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_5_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_6_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_7_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_8_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_9_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_10_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_11_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_12_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_13_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_14_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_15_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_16_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_17_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_18_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_19_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_20_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_21_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_22_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_23_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_24_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_25_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_26_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_27_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_28_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_29_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_30_owner; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_regStatus_31_owner; // @[Core_1.scala 88:23]
  wire  lsuRS_io_cdb_0_valid; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_cdb_0_bits_data; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_cdb_0_bits_id; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_cdb_0_bits_rd; // @[Core_1.scala 88:23]
  wire  lsuRS_io_cdb_1_valid; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_cdb_1_bits_data; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_cdb_1_bits_id; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_cdb_1_bits_rd; // @[Core_1.scala 88:23]
  wire  lsuRS_io_cdb_2_valid; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_cdb_2_bits_data; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_cdb_2_bits_id; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_cdb_2_bits_rd; // @[Core_1.scala 88:23]
  wire  lsuRS_io_cdb_3_valid; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_cdb_3_bits_data; // @[Core_1.scala 88:23]
  wire [7:0] lsuRS_io_cdb_3_bits_id; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_cdb_3_bits_rd; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_rf_0_addr; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_rf_0_data; // @[Core_1.scala 88:23]
  wire [4:0] lsuRS_io_rf_1_addr; // @[Core_1.scala 88:23]
  wire [31:0] lsuRS_io_rf_1_data; // @[Core_1.scala 88:23]
  wire  lsuRS_io_flush; // @[Core_1.scala 88:23]
  wire  csrStage_1_clock; // @[Core_1.scala 90:28]
  wire  csrStage_1_reset; // @[Core_1.scala 90:28]
  wire  csrStage_1_io_in_ready; // @[Core_1.scala 90:28]
  wire  csrStage_1_io_in_valid; // @[Core_1.scala 90:28]
  wire [2:0] csrStage_1_io_in_bits_csrOp; // @[Core_1.scala 90:28]
  wire [3:0] csrStage_1_io_in_bits_excpType; // @[Core_1.scala 90:28]
  wire [31:0] csrStage_1_io_in_bits_rs1Val; // @[Core_1.scala 90:28]
  wire [31:0] csrStage_1_io_in_bits_inst; // @[Core_1.scala 90:28]
  wire [7:0] csrStage_1_io_in_bits_id; // @[Core_1.scala 90:28]
  wire  csrStage_1_io_out_valid; // @[Core_1.scala 90:28]
  wire [4:0] csrStage_1_io_out_bits_rd; // @[Core_1.scala 90:28]
  wire [31:0] csrStage_1_io_out_bits_data; // @[Core_1.scala 90:28]
  wire [31:0] csrStage_1_io_out_bits_excpAddr; // @[Core_1.scala 90:28]
  wire  csrStage_1_io_out_bits_excpValid; // @[Core_1.scala 90:28]
  wire [7:0] csrStage_1_io_out_bits_id; // @[Core_1.scala 90:28]
  wire  csrStage_1_io_flush; // @[Core_1.scala 90:28]
  wire [31:0] csrStage_1_csrState_mcycle; // @[Core_1.scala 90:28]
  wire [31:0] csrStage_1_csrState_mcycleh; // @[Core_1.scala 90:28]
  wire  csrRS_clock; // @[Core_1.scala 91:23]
  wire  csrRS_reset; // @[Core_1.scala 91:23]
  wire  csrRS_io_enq_ready; // @[Core_1.scala 91:23]
  wire  csrRS_io_enq_valid; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_enq_bits_op; // @[Core_1.scala 91:23]
  wire [3:0] csrRS_io_enq_bits_opr1; // @[Core_1.scala 91:23]
  wire [3:0] csrRS_io_enq_bits_opr2; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_enq_bits_rs1; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_enq_bits_rs2; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_enq_bits_ROBId; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_enq_bits_rs1ROBId; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_enq_bits_rs2ROBId; // @[Core_1.scala 91:23]
  wire [2:0] csrRS_io_enq_bits_immSrc; // @[Core_1.scala 91:23]
  wire  csrRS_io_enq_bits_immSign; // @[Core_1.scala 91:23]
  wire [3:0] csrRS_io_enq_bits_excpType; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_enq_bits_pc; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_enq_bits_inst; // @[Core_1.scala 91:23]
  wire  csrRS_io_deq_ready; // @[Core_1.scala 91:23]
  wire  csrRS_io_deq_valid; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_deq_bits_op; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_deq_bits_ROBId; // @[Core_1.scala 91:23]
  wire [3:0] csrRS_io_deq_bits_opr1; // @[Core_1.scala 91:23]
  wire [3:0] csrRS_io_deq_bits_opr2; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_deq_bits_rs1Val; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_deq_bits_rs2Val; // @[Core_1.scala 91:23]
  wire [2:0] csrRS_io_deq_bits_immSrc; // @[Core_1.scala 91:23]
  wire  csrRS_io_deq_bits_immSign; // @[Core_1.scala 91:23]
  wire [3:0] csrRS_io_deq_bits_excpType; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_deq_bits_pc; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_deq_bits_inst; // @[Core_1.scala 91:23]
  wire  csrRS_io_robOut_valid; // @[Core_1.scala 91:23]
  wire [2:0] csrRS_io_robOut_bits_id; // @[Core_1.scala 91:23]
  wire  csrRS_io_robRead_0_busy; // @[Core_1.scala 91:23]
  wire [1:0] csrRS_io_robRead_0_state; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_robRead_0_rd; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_robRead_0_data; // @[Core_1.scala 91:23]
  wire  csrRS_io_robRead_1_busy; // @[Core_1.scala 91:23]
  wire [1:0] csrRS_io_robRead_1_state; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_robRead_1_rd; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_robRead_1_data; // @[Core_1.scala 91:23]
  wire  csrRS_io_robRead_2_busy; // @[Core_1.scala 91:23]
  wire [1:0] csrRS_io_robRead_2_state; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_robRead_2_rd; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_robRead_2_data; // @[Core_1.scala 91:23]
  wire  csrRS_io_robRead_3_busy; // @[Core_1.scala 91:23]
  wire [1:0] csrRS_io_robRead_3_state; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_robRead_3_rd; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_robRead_3_data; // @[Core_1.scala 91:23]
  wire  csrRS_io_robRead_4_busy; // @[Core_1.scala 91:23]
  wire [1:0] csrRS_io_robRead_4_state; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_robRead_4_rd; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_robRead_4_data; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_0_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_1_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_2_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_3_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_4_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_5_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_6_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_7_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_8_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_9_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_10_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_11_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_12_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_13_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_14_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_15_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_16_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_17_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_18_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_19_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_20_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_21_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_22_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_23_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_24_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_25_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_26_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_27_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_28_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_29_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_30_owner; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_regStatus_31_owner; // @[Core_1.scala 91:23]
  wire  csrRS_io_cdb_0_valid; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_cdb_0_bits_data; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_cdb_0_bits_id; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_cdb_0_bits_rd; // @[Core_1.scala 91:23]
  wire  csrRS_io_cdb_1_valid; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_cdb_1_bits_data; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_cdb_1_bits_id; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_cdb_1_bits_rd; // @[Core_1.scala 91:23]
  wire  csrRS_io_cdb_2_valid; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_cdb_2_bits_data; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_cdb_2_bits_id; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_cdb_2_bits_rd; // @[Core_1.scala 91:23]
  wire  csrRS_io_cdb_3_valid; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_cdb_3_bits_data; // @[Core_1.scala 91:23]
  wire [7:0] csrRS_io_cdb_3_bits_id; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_cdb_3_bits_rd; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_rf_0_addr; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_rf_0_data; // @[Core_1.scala 91:23]
  wire [4:0] csrRS_io_rf_1_addr; // @[Core_1.scala 91:23]
  wire [31:0] csrRS_io_rf_1_data; // @[Core_1.scala 91:23]
  wire  csrRS_io_flush; // @[Core_1.scala 91:23]
  wire  edgeBackPressure_clock; // @[Core_1.scala 130:34]
  wire  edgeBackPressure_io_in; // @[Core_1.scala 130:34]
  wire  edgeBackPressure_io_change; // @[Core_1.scala 130:34]
  wire  fetch_pendingBranch_clock; // @[Core_1.scala 135:37]
  wire  fetch_pendingBranch_reset; // @[Core_1.scala 135:37]
  wire  fetch_pendingBranch_io_enq_ready; // @[Core_1.scala 135:37]
  wire  fetch_pendingBranch_io_enq_valid; // @[Core_1.scala 135:37]
  wire [31:0] fetch_pendingBranch_io_enq_bits; // @[Core_1.scala 135:37]
  wire  fetch_pendingBranch_io_deq_ready; // @[Core_1.scala 135:37]
  wire  fetch_pendingBranch_io_deq_valid; // @[Core_1.scala 135:37]
  wire [31:0] fetch_pendingBranch_io_deq_bits; // @[Core_1.scala 135:37]
  wire [31:0] dec_decoders_0_io_inst; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_0_io_out_brType; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_0_io_out_wbType; // @[Core_1.scala 198:53]
  wire [4:0] dec_decoders_0_io_out_lsuOp; // @[Core_1.scala 198:53]
  wire [4:0] dec_decoders_0_io_out_aluOp; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_0_io_out_opr1; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_0_io_out_opr2; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_0_io_out_immSrc; // @[Core_1.scala 198:53]
  wire  dec_decoders_0_io_out_immSign; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_0_io_out_csrOp; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_0_io_out_excpType; // @[Core_1.scala 198:53]
  wire [31:0] dec_decoders_1_io_inst; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_1_io_out_brType; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_1_io_out_wbType; // @[Core_1.scala 198:53]
  wire [4:0] dec_decoders_1_io_out_lsuOp; // @[Core_1.scala 198:53]
  wire [4:0] dec_decoders_1_io_out_aluOp; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_1_io_out_opr1; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_1_io_out_opr2; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_1_io_out_immSrc; // @[Core_1.scala 198:53]
  wire  dec_decoders_1_io_out_immSign; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_1_io_out_csrOp; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_1_io_out_excpType; // @[Core_1.scala 198:53]
  wire [31:0] dec_decoders_2_io_inst; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_2_io_out_brType; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_2_io_out_wbType; // @[Core_1.scala 198:53]
  wire [4:0] dec_decoders_2_io_out_lsuOp; // @[Core_1.scala 198:53]
  wire [4:0] dec_decoders_2_io_out_aluOp; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_2_io_out_opr1; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_2_io_out_opr2; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_2_io_out_immSrc; // @[Core_1.scala 198:53]
  wire  dec_decoders_2_io_out_immSign; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_2_io_out_csrOp; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_2_io_out_excpType; // @[Core_1.scala 198:53]
  wire [31:0] dec_decoders_3_io_inst; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_3_io_out_brType; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_3_io_out_wbType; // @[Core_1.scala 198:53]
  wire [4:0] dec_decoders_3_io_out_lsuOp; // @[Core_1.scala 198:53]
  wire [4:0] dec_decoders_3_io_out_aluOp; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_3_io_out_opr1; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_3_io_out_opr2; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_3_io_out_immSrc; // @[Core_1.scala 198:53]
  wire  dec_decoders_3_io_out_immSign; // @[Core_1.scala 198:53]
  wire [2:0] dec_decoders_3_io_out_csrOp; // @[Core_1.scala 198:53]
  wire [3:0] dec_decoders_3_io_out_excpType; // @[Core_1.scala 198:53]
  wire  dcache_clock; // @[Core_1.scala 570:24]
  wire  dcache_reset; // @[Core_1.scala 570:24]
  wire  dcache_io_read_req_ready; // @[Core_1.scala 570:24]
  wire  dcache_io_read_req_valid; // @[Core_1.scala 570:24]
  wire [31:0] dcache_io_read_req_bits_addr; // @[Core_1.scala 570:24]
  wire  dcache_io_read_resp_ready; // @[Core_1.scala 570:24]
  wire  dcache_io_read_resp_valid; // @[Core_1.scala 570:24]
  wire [31:0] dcache_io_read_resp_bits_data; // @[Core_1.scala 570:24]
  wire  dcache_io_write_req_ready; // @[Core_1.scala 570:24]
  wire  dcache_io_write_req_valid; // @[Core_1.scala 570:24]
  wire [31:0] dcache_io_write_req_bits_addr; // @[Core_1.scala 570:24]
  wire [31:0] dcache_io_write_req_bits_data; // @[Core_1.scala 570:24]
  wire [3:0] dcache_io_write_req_bits_mask; // @[Core_1.scala 570:24]
  wire  dcache_io_write_resp_ready; // @[Core_1.scala 570:24]
  wire  dcache_io_write_resp_valid; // @[Core_1.scala 570:24]
  wire  dcache_io_tlbus_req_ready; // @[Core_1.scala 570:24]
  wire  dcache_io_tlbus_req_valid; // @[Core_1.scala 570:24]
  wire [2:0] dcache_io_tlbus_req_bits_opcode; // @[Core_1.scala 570:24]
  wire [31:0] dcache_io_tlbus_req_bits_address; // @[Core_1.scala 570:24]
  wire [127:0] dcache_io_tlbus_req_bits_data; // @[Core_1.scala 570:24]
  wire  dcache_io_tlbus_resp_valid; // @[Core_1.scala 570:24]
  wire [2:0] dcache_io_tlbus_resp_bits_opcode; // @[Core_1.scala 570:24]
  wire [127:0] dcache_io_tlbus_resp_bits_data; // @[Core_1.scala 570:24]
  wire  dcache_io_flush; // @[Core_1.scala 570:24]
  wire  xbar_clock; // @[Core_1.scala 695:22]
  wire  xbar_reset; // @[Core_1.scala 695:22]
  wire  xbar_io_masterFace_in_0_ready; // @[Core_1.scala 695:22]
  wire  xbar_io_masterFace_in_0_valid; // @[Core_1.scala 695:22]
  wire [31:0] xbar_io_masterFace_in_0_bits_address; // @[Core_1.scala 695:22]
  wire  xbar_io_masterFace_in_1_ready; // @[Core_1.scala 695:22]
  wire  xbar_io_masterFace_in_1_valid; // @[Core_1.scala 695:22]
  wire [2:0] xbar_io_masterFace_in_1_bits_opcode; // @[Core_1.scala 695:22]
  wire [31:0] xbar_io_masterFace_in_1_bits_address; // @[Core_1.scala 695:22]
  wire [127:0] xbar_io_masterFace_in_1_bits_data; // @[Core_1.scala 695:22]
  wire  xbar_io_masterFace_out_0_valid; // @[Core_1.scala 695:22]
  wire [2:0] xbar_io_masterFace_out_0_bits_opcode; // @[Core_1.scala 695:22]
  wire [127:0] xbar_io_masterFace_out_0_bits_data; // @[Core_1.scala 695:22]
  wire  xbar_io_masterFace_out_1_valid; // @[Core_1.scala 695:22]
  wire [2:0] xbar_io_masterFace_out_1_bits_opcode; // @[Core_1.scala 695:22]
  wire [127:0] xbar_io_masterFace_out_1_bits_data; // @[Core_1.scala 695:22]
  wire  xbar_io_slaveFace_in_0_ready; // @[Core_1.scala 695:22]
  wire  xbar_io_slaveFace_in_0_valid; // @[Core_1.scala 695:22]
  wire [2:0] xbar_io_slaveFace_in_0_bits_opcode; // @[Core_1.scala 695:22]
  wire [127:0] xbar_io_slaveFace_in_0_bits_size; // @[Core_1.scala 695:22]
  wire [31:0] xbar_io_slaveFace_in_0_bits_address; // @[Core_1.scala 695:22]
  wire [127:0] xbar_io_slaveFace_in_0_bits_data; // @[Core_1.scala 695:22]
  wire  xbar_io_slaveFace_out_0_ready; // @[Core_1.scala 695:22]
  wire  xbar_io_slaveFace_out_0_valid; // @[Core_1.scala 695:22]
  wire [2:0] xbar_io_slaveFace_out_0_bits_opcode; // @[Core_1.scala 695:22]
  wire [127:0] xbar_io_slaveFace_out_0_bits_data; // @[Core_1.scala 695:22]
  wire  rom_clock; // @[Core_1.scala 696:21]
  wire  rom_reset; // @[Core_1.scala 696:21]
  wire  rom_io_req_ready; // @[Core_1.scala 696:21]
  wire  rom_io_req_valid; // @[Core_1.scala 696:21]
  wire [2:0] rom_io_req_bits_opcode; // @[Core_1.scala 696:21]
  wire [127:0] rom_io_req_bits_size; // @[Core_1.scala 696:21]
  wire [31:0] rom_io_req_bits_address; // @[Core_1.scala 696:21]
  wire [127:0] rom_io_req_bits_data; // @[Core_1.scala 696:21]
  wire  rom_io_resp_ready; // @[Core_1.scala 696:21]
  wire  rom_io_resp_valid; // @[Core_1.scala 696:21]
  wire [2:0] rom_io_resp_bits_opcode; // @[Core_1.scala 696:21]
  wire [127:0] rom_io_resp_bits_size; // @[Core_1.scala 696:21]
  wire [127:0] rom_io_resp_bits_data; // @[Core_1.scala 696:21]
  wire  _csrExcpValid_T = rob_io_deq_ready & rob_io_deq_valid; // @[Decoupled.scala 51:35]
  wire  csrExcpValid = rob_io_deq_bits_excpValid & _csrExcpValid_T; // @[Core_1.scala 664:47]
  wire  bruBrTaken = rob_io_deq_bits_brTaken & _csrExcpValid_T; // @[Core_1.scala 662:43]
  wire  globalBrTaken = csrExcpValid | bruBrTaken; // @[Core_1.scala 104:38]
  wire [31:0] csrExcpAddr = rob_io_deq_bits_excpAddr; // @[Core_1.scala 102:31 665:17]
  wire [31:0] bruBrAddr = rob_io_deq_bits_brAddr; // @[Core_1.scala 663:15 99:29]
  wire [31:0] globalBrAddr = csrExcpValid ? csrExcpAddr : bruBrAddr; // @[Core_1.scala 105:27]
  reg [31:0] pcReg; // @[Core_1.scala 114:24]
  wire  isAlignAddr = ~(|pcReg[3:0]); // @[Core_1.scala 117:23]
  wire  _lastPc_T = icache_io_read_req_ready & icache_io_read_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] lastPc; // @[Reg.scala 19:16]
  wire [31:0] _pcNext4_T_1 = pcReg + 32'h10; // @[Core_1.scala 120:31]
  wire [4:0] _GEN_108 = {{1'd0}, lastPc[3:0]}; // @[Core_1.scala 121:45]
  wire [4:0] _pcNext4_T_4 = 5'h10 - _GEN_108; // @[Core_1.scala 121:45]
  wire [4:0] _pcNext4_T_6 = {_pcNext4_T_4[4:2], 2'h0}; // @[Core_1.scala 121:82]
  wire [31:0] _GEN_109 = {{27'd0}, _pcNext4_T_6}; // @[Core_1.scala 121:32]
  wire [31:0] _pcNext4_T_8 = lastPc + _GEN_109; // @[Core_1.scala 121:32]
  wire [31:0] pcNext4 = isAlignAddr ? _pcNext4_T_1 : _pcNext4_T_8; // @[Core_1.scala 119:22]
  reg  firstFire; // @[Reg.scala 35:20]
  wire  _GEN_3 = _lastPc_T ? 1'h0 : firstFire; // @[Reg.scala 36:18 35:20 36:22]
  wire  brTaken = fetch_pendingBranch_io_deq_ready & fetch_pendingBranch_io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _preFetchInst_T_2 = ~firstFire; // @[Core_1.scala 143:26]
  wire  fetch_fire = icache_io_read_resp_valid; // @[Core_1.scala 161:17 94:27]
  wire  _preFetchInst_T_6 = (fetch_fire | edgeBackPressure_io_change) & ~ib_io_status_back_pressure | brTaken; // @[Core_1.scala 144:107]
  wire  _preFetchInst_T_7 = ~firstFire & _preFetchInst_T_6; // @[Core_1.scala 143:37]
  wire  preFetchInst = firstFire & pcReg == 32'h0 | _preFetchInst_T_7; // @[Core_1.scala 142:59]
  wire [31:0] pcNext = brTaken ? fetch_pendingBranch_io_deq_bits : pcNext4; // @[Core_1.scala 159:18]
  wire [31:0] _icache_io_read_req_bits_addr_T_1 = firstFire ? pcReg : pcNext; // @[Core_1.scala 151:69]
  wire [31:0] _icache_io_read_req_bits_addr_T_2 = brTaken ? fetch_pendingBranch_io_deq_bits : pcReg; // @[Core_1.scala 151:100]
  reg [31:0] blockAddr; // @[Reg.scala 19:16]
  reg  blockValid; // @[Core_1.scala 166:29]
  wire  willBlock = (globalBrTaken | brTaken) & icache_io_read_resp_bits_addr != globalBrAddr; // @[Core_1.scala 167:48]
  wire  willWakeUp = blockValid & icache_io_read_resp_valid & icache_io_read_resp_bits_addr == blockAddr; // @[Core_1.scala 168:62]
  wire  _GEN_6 = willWakeUp ? 1'h0 : blockValid; // @[Core_1.scala 170:27 166:29 170:40]
  wire  _GEN_7 = willBlock | _GEN_6; // @[Core_1.scala 169:{21,34}]
  wire  icacheRespIsAlignAddr = ~(|icache_io_read_resp_bits_addr[3:0]); // @[Core_1.scala 109:9]
  wire [2:0] _GEN_110 = {{1'd0}, icache_io_read_resp_bits_addr[3:2]}; // @[Core_1.scala 177:93]
  wire [2:0] _ib_io_in_bits_icache_size_T_2 = 3'h4 - _GEN_110; // @[Core_1.scala 177:93]
  wire  _ib_io_in_bits_flush_T_1 = globalBrTaken | reset; // @[Core_1.scala 179:42]
  reg  dec_full; // @[Core_1.scala 186:27]
  wire  _dec_valid_T = ~_ib_io_in_bits_flush_T_1; // @[Core_1.scala 209:30]
  wire  dec_valid = dec_full & ~_ib_io_in_bits_flush_T_1; // @[Core_1.scala 209:27]
  reg  issue_full; // @[Core_1.scala 224:29]
  wire  _issue_ready_T = ~issue_full; // @[Core_1.scala 241:20]
  reg [1:0] issue_ptr; // @[Core_1.scala 231:28]
  reg [3:0] issue_instValid; // @[Reg.scala 19:16]
  wire [1:0] _issue_instSize_T_4 = issue_instValid[0] + issue_instValid[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _issue_instSize_T_6 = issue_instValid[2] + issue_instValid[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _issue_instSize_T_8 = _issue_instSize_T_4 + _issue_instSize_T_6; // @[Bitwise.scala 51:90]
  wire [2:0] issue_instSize = _issue_instSize_T_8 - 3'h1; // @[Core_1.scala 229:52]
  wire [2:0] _GEN_111 = {{1'd0}, issue_ptr}; // @[Core_1.scala 247:32]
  wire  issue_instFire = rob_io_enq_ready & rob_io_enq_valid; // @[Decoupled.scala 51:35]
  wire  issue_fire = _GEN_111 == issue_instSize & issue_instFire & _dec_valid_T; // @[Core_1.scala 247:71]
  wire  issue_ready = ~issue_full | issue_fire; // @[Core_1.scala 241:32]
  wire  dec_fire = dec_valid & issue_ready; // @[Core_1.scala 187:30]
  wire  dec_ready = ~dec_full | dec_fire; // @[Core_1.scala 193:28]
  wire  dec_latch = ib_io_out_valid & dec_ready; // @[Core_1.scala 185:37]
  reg [31:0] dec_inst_0_inst; // @[Reg.scala 19:16]
  reg  dec_inst_0_valid; // @[Reg.scala 19:16]
  reg [31:0] dec_inst_1_inst; // @[Reg.scala 19:16]
  reg  dec_inst_1_valid; // @[Reg.scala 19:16]
  reg [31:0] dec_inst_2_inst; // @[Reg.scala 19:16]
  reg  dec_inst_2_valid; // @[Reg.scala 19:16]
  reg [31:0] dec_inst_3_inst; // @[Reg.scala 19:16]
  reg  dec_inst_3_valid; // @[Reg.scala 19:16]
  reg [31:0] dec_pc; // @[Reg.scala 19:16]
  wire  _GEN_17 = dec_full & dec_fire ? 1'h0 : dec_full; // @[Core_1.scala 186:27 195:{37,48}]
  wire  _GEN_18 = dec_latch | _GEN_17; // @[Core_1.scala 194:{21,32}]
  reg [31:0] issue_pc; // @[Reg.scala 19:16]
  reg [3:0] issue_decodeSigs_0_brType; // @[Core_1.scala 226:31]
  reg [4:0] issue_decodeSigs_0_lsuOp; // @[Core_1.scala 226:31]
  reg [4:0] issue_decodeSigs_0_aluOp; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_0_opr1; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_0_opr2; // @[Core_1.scala 226:31]
  reg [2:0] issue_decodeSigs_0_immSrc; // @[Core_1.scala 226:31]
  reg  issue_decodeSigs_0_immSign; // @[Core_1.scala 226:31]
  reg [2:0] issue_decodeSigs_0_csrOp; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_0_excpType; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_1_brType; // @[Core_1.scala 226:31]
  reg [4:0] issue_decodeSigs_1_lsuOp; // @[Core_1.scala 226:31]
  reg [4:0] issue_decodeSigs_1_aluOp; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_1_opr1; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_1_opr2; // @[Core_1.scala 226:31]
  reg [2:0] issue_decodeSigs_1_immSrc; // @[Core_1.scala 226:31]
  reg  issue_decodeSigs_1_immSign; // @[Core_1.scala 226:31]
  reg [2:0] issue_decodeSigs_1_csrOp; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_1_excpType; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_2_brType; // @[Core_1.scala 226:31]
  reg [4:0] issue_decodeSigs_2_lsuOp; // @[Core_1.scala 226:31]
  reg [4:0] issue_decodeSigs_2_aluOp; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_2_opr1; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_2_opr2; // @[Core_1.scala 226:31]
  reg [2:0] issue_decodeSigs_2_immSrc; // @[Core_1.scala 226:31]
  reg  issue_decodeSigs_2_immSign; // @[Core_1.scala 226:31]
  reg [2:0] issue_decodeSigs_2_csrOp; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_2_excpType; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_3_brType; // @[Core_1.scala 226:31]
  reg [4:0] issue_decodeSigs_3_lsuOp; // @[Core_1.scala 226:31]
  reg [4:0] issue_decodeSigs_3_aluOp; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_3_opr1; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_3_opr2; // @[Core_1.scala 226:31]
  reg [2:0] issue_decodeSigs_3_immSrc; // @[Core_1.scala 226:31]
  reg  issue_decodeSigs_3_immSign; // @[Core_1.scala 226:31]
  reg [2:0] issue_decodeSigs_3_csrOp; // @[Core_1.scala 226:31]
  reg [3:0] issue_decodeSigs_3_excpType; // @[Core_1.scala 226:31]
  wire [3:0] _issue_instValid_T = {dec_inst_0_valid,dec_inst_1_valid,dec_inst_2_valid,dec_inst_3_valid}; // @[Cat.scala 33:92]
  reg [31:0] issue_inst_0; // @[Core_1.scala 228:25]
  reg [31:0] issue_inst_1; // @[Core_1.scala 228:25]
  reg [31:0] issue_inst_2; // @[Core_1.scala 228:25]
  reg [31:0] issue_inst_3; // @[Core_1.scala 228:25]
  wire [3:0] dec_decodeSigs_0_brType = dec_decoders_0_io_out_brType; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_0_wbType = dec_decoders_0_io_out_wbType; // @[Core_1.scala 199:57 202:27]
  wire [4:0] dec_decodeSigs_0_lsuOp = dec_decoders_0_io_out_lsuOp; // @[Core_1.scala 199:57 202:27]
  wire [4:0] dec_decodeSigs_0_aluOp = dec_decoders_0_io_out_aluOp; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_0_opr1 = dec_decoders_0_io_out_opr1; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_0_opr2 = dec_decoders_0_io_out_opr2; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_0_immSrc = dec_decoders_0_io_out_immSrc; // @[Core_1.scala 199:57 202:27]
  wire  dec_decodeSigs_0_immSign = dec_decoders_0_io_out_immSign; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_0_csrOp = dec_decoders_0_io_out_csrOp; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_0_excpType = dec_decoders_0_io_out_excpType; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_1_brType = dec_decoders_1_io_out_brType; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_1_wbType = dec_decoders_1_io_out_wbType; // @[Core_1.scala 199:57 202:27]
  wire [4:0] dec_decodeSigs_1_lsuOp = dec_decoders_1_io_out_lsuOp; // @[Core_1.scala 199:57 202:27]
  wire [4:0] dec_decodeSigs_1_aluOp = dec_decoders_1_io_out_aluOp; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_1_opr1 = dec_decoders_1_io_out_opr1; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_1_opr2 = dec_decoders_1_io_out_opr2; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_1_immSrc = dec_decoders_1_io_out_immSrc; // @[Core_1.scala 199:57 202:27]
  wire  dec_decodeSigs_1_immSign = dec_decoders_1_io_out_immSign; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_1_csrOp = dec_decoders_1_io_out_csrOp; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_1_excpType = dec_decoders_1_io_out_excpType; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_2_brType = dec_decoders_2_io_out_brType; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_2_wbType = dec_decoders_2_io_out_wbType; // @[Core_1.scala 199:57 202:27]
  wire [4:0] dec_decodeSigs_2_lsuOp = dec_decoders_2_io_out_lsuOp; // @[Core_1.scala 199:57 202:27]
  wire [4:0] dec_decodeSigs_2_aluOp = dec_decoders_2_io_out_aluOp; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_2_opr1 = dec_decoders_2_io_out_opr1; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_2_opr2 = dec_decoders_2_io_out_opr2; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_2_immSrc = dec_decoders_2_io_out_immSrc; // @[Core_1.scala 199:57 202:27]
  wire  dec_decodeSigs_2_immSign = dec_decoders_2_io_out_immSign; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_2_csrOp = dec_decoders_2_io_out_csrOp; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_2_excpType = dec_decoders_2_io_out_excpType; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_3_brType = dec_decoders_3_io_out_brType; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_3_wbType = dec_decoders_3_io_out_wbType; // @[Core_1.scala 199:57 202:27]
  wire [4:0] dec_decodeSigs_3_lsuOp = dec_decoders_3_io_out_lsuOp; // @[Core_1.scala 199:57 202:27]
  wire [4:0] dec_decodeSigs_3_aluOp = dec_decoders_3_io_out_aluOp; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_3_opr1 = dec_decoders_3_io_out_opr1; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_3_opr2 = dec_decoders_3_io_out_opr2; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_3_immSrc = dec_decoders_3_io_out_immSrc; // @[Core_1.scala 199:57 202:27]
  wire  dec_decodeSigs_3_immSign = dec_decoders_3_io_out_immSign; // @[Core_1.scala 199:57 202:27]
  wire [2:0] dec_decodeSigs_3_csrOp = dec_decoders_3_io_out_csrOp; // @[Core_1.scala 199:57 202:27]
  wire [3:0] dec_decodeSigs_3_excpType = dec_decoders_3_io_out_excpType; // @[Core_1.scala 199:57 202:27]
  wire  _GEN_70 = issue_full & issue_fire ? 1'h0 : issue_full; // @[Core_1.scala 224:29 243:{41,54}]
  wire  _GEN_71 = dec_fire | _GEN_70; // @[Core_1.scala 242:{23,36}]
  wire [1:0] _issue_ptr_T_1 = issue_ptr + 2'h1; // @[Core_1.scala 249:56]
  wire [3:0] _issue_chosenDecodesigs_T = 4'h1 << issue_ptr; // @[OneHot.scala 57:35]
  wire [3:0] _issue_chosenDecodesigs_T_5 = _issue_chosenDecodesigs_T[0] ? issue_decodeSigs_0_excpType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_6 = _issue_chosenDecodesigs_T[1] ? issue_decodeSigs_1_excpType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_7 = _issue_chosenDecodesigs_T[2] ? issue_decodeSigs_2_excpType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_8 = _issue_chosenDecodesigs_T[3] ? issue_decodeSigs_3_excpType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_9 = _issue_chosenDecodesigs_T_5 | _issue_chosenDecodesigs_T_6; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_10 = _issue_chosenDecodesigs_T_9 | _issue_chosenDecodesigs_T_7; // @[Mux.scala 27:73]
  wire [3:0] issue_chosenDecodesigs_excpType = _issue_chosenDecodesigs_T_10 | _issue_chosenDecodesigs_T_8; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_12 = _issue_chosenDecodesigs_T[0] ? issue_decodeSigs_0_csrOp : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_13 = _issue_chosenDecodesigs_T[1] ? issue_decodeSigs_1_csrOp : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_14 = _issue_chosenDecodesigs_T[2] ? issue_decodeSigs_2_csrOp : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_15 = _issue_chosenDecodesigs_T[3] ? issue_decodeSigs_3_csrOp : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_16 = _issue_chosenDecodesigs_T_12 | _issue_chosenDecodesigs_T_13; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_17 = _issue_chosenDecodesigs_T_16 | _issue_chosenDecodesigs_T_14; // @[Mux.scala 27:73]
  wire [2:0] issue_chosenDecodesigs_csrOp = _issue_chosenDecodesigs_T_17 | _issue_chosenDecodesigs_T_15; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_26 = _issue_chosenDecodesigs_T[0] ? issue_decodeSigs_0_immSrc : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_27 = _issue_chosenDecodesigs_T[1] ? issue_decodeSigs_1_immSrc : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_28 = _issue_chosenDecodesigs_T[2] ? issue_decodeSigs_2_immSrc : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_29 = _issue_chosenDecodesigs_T[3] ? issue_decodeSigs_3_immSrc : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_30 = _issue_chosenDecodesigs_T_26 | _issue_chosenDecodesigs_T_27; // @[Mux.scala 27:73]
  wire [2:0] _issue_chosenDecodesigs_T_31 = _issue_chosenDecodesigs_T_30 | _issue_chosenDecodesigs_T_28; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_33 = _issue_chosenDecodesigs_T[0] ? issue_decodeSigs_0_opr2 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_34 = _issue_chosenDecodesigs_T[1] ? issue_decodeSigs_1_opr2 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_35 = _issue_chosenDecodesigs_T[2] ? issue_decodeSigs_2_opr2 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_36 = _issue_chosenDecodesigs_T[3] ? issue_decodeSigs_3_opr2 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_37 = _issue_chosenDecodesigs_T_33 | _issue_chosenDecodesigs_T_34; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_38 = _issue_chosenDecodesigs_T_37 | _issue_chosenDecodesigs_T_35; // @[Mux.scala 27:73]
  wire [3:0] issue_chosenDecodesigs_opr2 = _issue_chosenDecodesigs_T_38 | _issue_chosenDecodesigs_T_36; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_40 = _issue_chosenDecodesigs_T[0] ? issue_decodeSigs_0_opr1 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_41 = _issue_chosenDecodesigs_T[1] ? issue_decodeSigs_1_opr1 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_42 = _issue_chosenDecodesigs_T[2] ? issue_decodeSigs_2_opr1 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_43 = _issue_chosenDecodesigs_T[3] ? issue_decodeSigs_3_opr1 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_44 = _issue_chosenDecodesigs_T_40 | _issue_chosenDecodesigs_T_41; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_45 = _issue_chosenDecodesigs_T_44 | _issue_chosenDecodesigs_T_42; // @[Mux.scala 27:73]
  wire [3:0] issue_chosenDecodesigs_opr1 = _issue_chosenDecodesigs_T_45 | _issue_chosenDecodesigs_T_43; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_47 = _issue_chosenDecodesigs_T[0] ? issue_decodeSigs_0_aluOp : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_48 = _issue_chosenDecodesigs_T[1] ? issue_decodeSigs_1_aluOp : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_49 = _issue_chosenDecodesigs_T[2] ? issue_decodeSigs_2_aluOp : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_50 = _issue_chosenDecodesigs_T[3] ? issue_decodeSigs_3_aluOp : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_51 = _issue_chosenDecodesigs_T_47 | _issue_chosenDecodesigs_T_48; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_52 = _issue_chosenDecodesigs_T_51 | _issue_chosenDecodesigs_T_49; // @[Mux.scala 27:73]
  wire [4:0] issue_chosenDecodesigs_aluOp = _issue_chosenDecodesigs_T_52 | _issue_chosenDecodesigs_T_50; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_54 = _issue_chosenDecodesigs_T[0] ? issue_decodeSigs_0_lsuOp : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_55 = _issue_chosenDecodesigs_T[1] ? issue_decodeSigs_1_lsuOp : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_56 = _issue_chosenDecodesigs_T[2] ? issue_decodeSigs_2_lsuOp : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_57 = _issue_chosenDecodesigs_T[3] ? issue_decodeSigs_3_lsuOp : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_58 = _issue_chosenDecodesigs_T_54 | _issue_chosenDecodesigs_T_55; // @[Mux.scala 27:73]
  wire [4:0] _issue_chosenDecodesigs_T_59 = _issue_chosenDecodesigs_T_58 | _issue_chosenDecodesigs_T_56; // @[Mux.scala 27:73]
  wire [4:0] issue_chosenDecodesigs_lsuOp = _issue_chosenDecodesigs_T_59 | _issue_chosenDecodesigs_T_57; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_68 = _issue_chosenDecodesigs_T[0] ? issue_decodeSigs_0_brType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_69 = _issue_chosenDecodesigs_T[1] ? issue_decodeSigs_1_brType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_70 = _issue_chosenDecodesigs_T[2] ? issue_decodeSigs_2_brType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_71 = _issue_chosenDecodesigs_T[3] ? issue_decodeSigs_3_brType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_72 = _issue_chosenDecodesigs_T_68 | _issue_chosenDecodesigs_T_69; // @[Mux.scala 27:73]
  wire [3:0] _issue_chosenDecodesigs_T_73 = _issue_chosenDecodesigs_T_72 | _issue_chosenDecodesigs_T_70; // @[Mux.scala 27:73]
  wire [3:0] issue_chosenDecodesigs_brType = _issue_chosenDecodesigs_T_73 | _issue_chosenDecodesigs_T_71; // @[Mux.scala 27:73]
  wire [31:0] _issue_chosenInst_T_5 = _issue_chosenDecodesigs_T[0] ? issue_inst_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _issue_chosenInst_T_6 = _issue_chosenDecodesigs_T[1] ? issue_inst_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _issue_chosenInst_T_7 = _issue_chosenDecodesigs_T[2] ? issue_inst_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _issue_chosenInst_T_8 = _issue_chosenDecodesigs_T[3] ? issue_inst_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _issue_chosenInst_T_9 = _issue_chosenInst_T_5 | _issue_chosenInst_T_6; // @[Mux.scala 27:73]
  wire [31:0] _issue_chosenInst_T_10 = _issue_chosenInst_T_9 | _issue_chosenInst_T_7; // @[Mux.scala 27:73]
  wire [31:0] issue_chosenInst = _issue_chosenInst_T_10 | _issue_chosenInst_T_8; // @[Mux.scala 27:73]
  wire [4:0] rs1 = issue_chosenInst[19:15]; // @[util.scala 72:31]
  wire [4:0] rs2 = issue_chosenInst[24:20]; // @[util.scala 73:31]
  wire [4:0] issue_rs1 = issue_chosenDecodesigs_opr1 == 4'h1 ? rs1 : 5'h0; // @[Core_1.scala 266:24]
  wire  issue_aluValid = issue_chosenDecodesigs_aluOp != 5'h11 & issue_full; // @[Core_1.scala 272:67]
  wire  issue_bruValid = issue_chosenDecodesigs_brType != 4'h0 & issue_full; // @[Core_1.scala 273:67]
  wire  issue_lsuValid = issue_chosenDecodesigs_lsuOp != 5'h0 & issue_full; // @[Core_1.scala 274:67]
  wire  issue_csrValid = (issue_chosenDecodesigs_csrOp != 3'h0 | issue_chosenDecodesigs_excpType != 4'h0) & issue_full; // @[Core_1.scala 275:117]
  wire [1:0] _T_8 = issue_aluValid + issue_bruValid; // @[Bitwise.scala 51:90]
  wire [1:0] _T_10 = issue_lsuValid + issue_csrValid; // @[Bitwise.scala 51:90]
  wire [2:0] _T_12 = _T_8 + _T_10; // @[Bitwise.scala 51:90]
  wire [3:0] _issue_stagePc_T = {issue_ptr, 2'h0}; // @[Core_1.scala 319:47]
  wire [31:0] _GEN_112 = {{28'd0}, _issue_stagePc_T}; // @[Core_1.scala 319:34]
  wire [31:0] issue_stagePc = issue_pc + _GEN_112; // @[Core_1.scala 319:34]
  wire  _rsReady_T_1 = issue_lsuValid ? lsuRS_io_enq_ready : issue_csrValid & csrRS_io_enq_ready; // @[Mux.scala 101:16]
  wire  _rsReady_T_2 = issue_bruValid ? bruRS_io_enq_ready : _rsReady_T_1; // @[Mux.scala 101:16]
  wire  rsReady = issue_aluValid ? aluRS_io_enq_ready : _rsReady_T_2; // @[Mux.scala 101:16]
  wire [4:0] _rob_io_enq_bits_fuOp_T = issue_csrValid ? {{2'd0}, issue_chosenDecodesigs_csrOp} : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _rob_io_enq_bits_fuOp_T_1 = issue_lsuValid ? issue_chosenDecodesigs_lsuOp : _rob_io_enq_bits_fuOp_T; // @[Mux.scala 101:16]
  wire [4:0] _rob_io_enq_bits_fuOp_T_2 = issue_bruValid ? {{1'd0}, issue_chosenDecodesigs_brType} :
    _rob_io_enq_bits_fuOp_T_1; // @[Mux.scala 101:16]
  wire [4:0] _rob_io_enq_bits_fuOp_T_3 = issue_aluValid ? issue_chosenDecodesigs_aluOp : _rob_io_enq_bits_fuOp_T_2; // @[Mux.scala 101:16]
  wire [1:0] rob_io_enq_bits_fuValid_lo = {issue_bruValid,issue_aluValid}; // @[Cat.scala 33:92]
  wire [1:0] rob_io_enq_bits_fuValid_hi = {issue_csrValid,issue_lsuValid}; // @[Cat.scala 33:92]
  wire [4:0] rd = issue_chosenInst[11:7]; // @[util.scala 71:31]
  wire [3:0] _invalidBRU_T = {{1'd0}, rob_io_enq_bits_fuValid[3:1]}; // @[Core_1.scala 474:33]
  wire  invalidBRU = _invalidBRU_T[0] & (rob_io_enq_bits_fuOp != 8'h2 & rob_io_enq_bits_fuOp != 8'h1); // @[Core_1.scala 474:39]
  wire [3:0] _invalidLSU_T = {{2'd0}, rob_io_enq_bits_fuValid[3:2]}; // @[Core_1.scala 475:33]
  wire  invalidLSU = _invalidLSU_T[0] & (rob_io_enq_bits_fuOp == 8'h8 | rob_io_enq_bits_fuOp == 8'h7 |
    rob_io_enq_bits_fuOp == 8'h6 | rob_io_enq_bits_fuOp == 8'h14); // @[Core_1.scala 475:39]
  wire  invalidRd = invalidBRU | invalidLSU | rd == 5'h0; // @[Core_1.scala 476:46]
  wire [7:0] _GEN_76 = rob_io_regStatus_0_owner; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_77 = 5'h1 == issue_rs1 ? rob_io_regStatus_1_owner : _GEN_76; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_78 = 5'h2 == issue_rs1 ? rob_io_regStatus_2_owner : _GEN_77; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_79 = 5'h3 == issue_rs1 ? rob_io_regStatus_3_owner : _GEN_78; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_80 = 5'h4 == issue_rs1 ? rob_io_regStatus_4_owner : _GEN_79; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_81 = 5'h5 == issue_rs1 ? rob_io_regStatus_5_owner : _GEN_80; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_82 = 5'h6 == issue_rs1 ? rob_io_regStatus_6_owner : _GEN_81; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_83 = 5'h7 == issue_rs1 ? rob_io_regStatus_7_owner : _GEN_82; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_84 = 5'h8 == issue_rs1 ? rob_io_regStatus_8_owner : _GEN_83; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_85 = 5'h9 == issue_rs1 ? rob_io_regStatus_9_owner : _GEN_84; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_86 = 5'ha == issue_rs1 ? rob_io_regStatus_10_owner : _GEN_85; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_87 = 5'hb == issue_rs1 ? rob_io_regStatus_11_owner : _GEN_86; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_88 = 5'hc == issue_rs1 ? rob_io_regStatus_12_owner : _GEN_87; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_89 = 5'hd == issue_rs1 ? rob_io_regStatus_13_owner : _GEN_88; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_90 = 5'he == issue_rs1 ? rob_io_regStatus_14_owner : _GEN_89; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_91 = 5'hf == issue_rs1 ? rob_io_regStatus_15_owner : _GEN_90; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_92 = 5'h10 == issue_rs1 ? rob_io_regStatus_16_owner : _GEN_91; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_93 = 5'h11 == issue_rs1 ? rob_io_regStatus_17_owner : _GEN_92; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_94 = 5'h12 == issue_rs1 ? rob_io_regStatus_18_owner : _GEN_93; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_95 = 5'h13 == issue_rs1 ? rob_io_regStatus_19_owner : _GEN_94; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_96 = 5'h14 == issue_rs1 ? rob_io_regStatus_20_owner : _GEN_95; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_97 = 5'h15 == issue_rs1 ? rob_io_regStatus_21_owner : _GEN_96; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_98 = 5'h16 == issue_rs1 ? rob_io_regStatus_22_owner : _GEN_97; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_99 = 5'h17 == issue_rs1 ? rob_io_regStatus_23_owner : _GEN_98; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_100 = 5'h18 == issue_rs1 ? rob_io_regStatus_24_owner : _GEN_99; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_101 = 5'h19 == issue_rs1 ? rob_io_regStatus_25_owner : _GEN_100; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_102 = 5'h1a == issue_rs1 ? rob_io_regStatus_26_owner : _GEN_101; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_103 = 5'h1b == issue_rs1 ? rob_io_regStatus_27_owner : _GEN_102; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_104 = 5'h1c == issue_rs1 ? rob_io_regStatus_28_owner : _GEN_103; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_105 = 5'h1d == issue_rs1 ? rob_io_regStatus_29_owner : _GEN_104; // @[Core_1.scala 500:{22,22}]
  wire [7:0] _GEN_106 = 5'h1e == issue_rs1 ? rob_io_regStatus_30_owner : _GEN_105; // @[Core_1.scala 500:{22,22}]
  reg  io_out_state_instState_REG_commit; // @[Core_1.scala 687:38]
  reg [31:0] io_out_state_instState_REG_pc; // @[Core_1.scala 687:38]
  reg [31:0] io_out_state_instState_REG_inst; // @[Core_1.scala 687:38]
  InstBuffer ib ( // @[Core_1.scala 50:20]
    .clock(ib_clock),
    .reset(ib_reset),
    .io_in_ready(ib_io_in_ready),
    .io_in_valid(ib_io_in_valid),
    .io_in_bits_icache_data(ib_io_in_bits_icache_data),
    .io_in_bits_icache_addr(ib_io_in_bits_icache_addr),
    .io_in_bits_icache_inst_0(ib_io_in_bits_icache_inst_0),
    .io_in_bits_icache_inst_1(ib_io_in_bits_icache_inst_1),
    .io_in_bits_icache_inst_2(ib_io_in_bits_icache_inst_2),
    .io_in_bits_icache_inst_3(ib_io_in_bits_icache_inst_3),
    .io_in_bits_icache_size(ib_io_in_bits_icache_size),
    .io_in_bits_pc(ib_io_in_bits_pc),
    .io_in_bits_flush(ib_io_in_bits_flush),
    .io_out_ready(ib_io_out_ready),
    .io_out_valid(ib_io_out_valid),
    .io_out_bits_inst_0_inst(ib_io_out_bits_inst_0_inst),
    .io_out_bits_inst_0_valid(ib_io_out_bits_inst_0_valid),
    .io_out_bits_inst_1_inst(ib_io_out_bits_inst_1_inst),
    .io_out_bits_inst_1_valid(ib_io_out_bits_inst_1_valid),
    .io_out_bits_inst_2_inst(ib_io_out_bits_inst_2_inst),
    .io_out_bits_inst_2_valid(ib_io_out_bits_inst_2_valid),
    .io_out_bits_inst_3_inst(ib_io_out_bits_inst_3_inst),
    .io_out_bits_inst_3_valid(ib_io_out_bits_inst_3_valid),
    .io_out_bits_pc(ib_io_out_bits_pc),
    .io_status_back_pressure(ib_io_status_back_pressure),
    .io_status_full(ib_io_status_full)
  );
  ICache icache ( // @[Core_1.scala 52:24]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_read_req_ready(icache_io_read_req_ready),
    .io_read_req_valid(icache_io_read_req_valid),
    .io_read_req_bits_addr(icache_io_read_req_bits_addr),
    .io_read_resp_ready(icache_io_read_resp_ready),
    .io_read_resp_valid(icache_io_read_resp_valid),
    .io_read_resp_bits_data(icache_io_read_resp_bits_data),
    .io_read_resp_bits_addr(icache_io_read_resp_bits_addr),
    .io_read_resp_bits_inst_0(icache_io_read_resp_bits_inst_0),
    .io_read_resp_bits_inst_1(icache_io_read_resp_bits_inst_1),
    .io_read_resp_bits_inst_2(icache_io_read_resp_bits_inst_2),
    .io_read_resp_bits_inst_3(icache_io_read_resp_bits_inst_3),
    .io_read_resp_bits_size(icache_io_read_resp_bits_size),
    .io_tlbus_req_ready(icache_io_tlbus_req_ready),
    .io_tlbus_req_valid(icache_io_tlbus_req_valid),
    .io_tlbus_req_bits_address(icache_io_tlbus_req_bits_address),
    .io_tlbus_resp_ready(icache_io_tlbus_resp_ready),
    .io_tlbus_resp_valid(icache_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(icache_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(icache_io_tlbus_resp_bits_data),
    .io_flush(icache_io_flush)
  );
  RegFile2 rf ( // @[Core_1.scala 64:20]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_r_0_addr(rf_io_r_0_addr),
    .io_r_0_data(rf_io_r_0_data),
    .io_r_1_addr(rf_io_r_1_addr),
    .io_r_1_data(rf_io_r_1_data),
    .io_r_2_addr(rf_io_r_2_addr),
    .io_r_2_data(rf_io_r_2_data),
    .io_r_3_addr(rf_io_r_3_addr),
    .io_r_3_data(rf_io_r_3_data),
    .io_r_4_addr(rf_io_r_4_addr),
    .io_r_4_data(rf_io_r_4_data),
    .io_r_5_addr(rf_io_r_5_addr),
    .io_r_5_data(rf_io_r_5_data),
    .io_r_6_addr(rf_io_r_6_addr),
    .io_r_6_data(rf_io_r_6_data),
    .io_r_7_addr(rf_io_r_7_addr),
    .io_r_7_data(rf_io_r_7_data),
    .io_w_0_addr(rf_io_w_0_addr),
    .io_w_0_en(rf_io_w_0_en),
    .io_w_0_data(rf_io_w_0_data),
    .regState_0_regState_0(rf_regState_0_regState_0),
    .regState_0_regState_1(rf_regState_0_regState_1),
    .regState_0_regState_2(rf_regState_0_regState_2),
    .regState_0_regState_3(rf_regState_0_regState_3),
    .regState_0_regState_4(rf_regState_0_regState_4),
    .regState_0_regState_5(rf_regState_0_regState_5),
    .regState_0_regState_6(rf_regState_0_regState_6),
    .regState_0_regState_7(rf_regState_0_regState_7),
    .regState_0_regState_8(rf_regState_0_regState_8),
    .regState_0_regState_9(rf_regState_0_regState_9),
    .regState_0_regState_10(rf_regState_0_regState_10),
    .regState_0_regState_11(rf_regState_0_regState_11),
    .regState_0_regState_12(rf_regState_0_regState_12),
    .regState_0_regState_13(rf_regState_0_regState_13),
    .regState_0_regState_14(rf_regState_0_regState_14),
    .regState_0_regState_15(rf_regState_0_regState_15),
    .regState_0_regState_16(rf_regState_0_regState_16),
    .regState_0_regState_17(rf_regState_0_regState_17),
    .regState_0_regState_18(rf_regState_0_regState_18),
    .regState_0_regState_19(rf_regState_0_regState_19),
    .regState_0_regState_20(rf_regState_0_regState_20),
    .regState_0_regState_21(rf_regState_0_regState_21),
    .regState_0_regState_22(rf_regState_0_regState_22),
    .regState_0_regState_23(rf_regState_0_regState_23),
    .regState_0_regState_24(rf_regState_0_regState_24),
    .regState_0_regState_25(rf_regState_0_regState_25),
    .regState_0_regState_26(rf_regState_0_regState_26),
    .regState_0_regState_27(rf_regState_0_regState_27),
    .regState_0_regState_28(rf_regState_0_regState_28),
    .regState_0_regState_29(rf_regState_0_regState_29),
    .regState_0_regState_30(rf_regState_0_regState_30),
    .regState_0_regState_31(rf_regState_0_regState_31)
  );
  ROB rob ( // @[Core_1.scala 79:21]
    .clock(rob_clock),
    .reset(rob_reset),
    .io_enq_ready(rob_io_enq_ready),
    .io_enq_valid(rob_io_enq_valid),
    .io_enq_bits_rd(rob_io_enq_bits_rd),
    .io_enq_bits_fuValid(rob_io_enq_bits_fuValid),
    .io_enq_bits_fuOp(rob_io_enq_bits_fuOp),
    .io_enq_bits_pc(rob_io_enq_bits_pc),
    .io_enq_bits_inst(rob_io_enq_bits_inst),
    .io_deq_ready(rob_io_deq_ready),
    .io_deq_valid(rob_io_deq_valid),
    .io_deq_bits_rdWrEn(rob_io_deq_bits_rdWrEn),
    .io_deq_bits_rd(rob_io_deq_bits_rd),
    .io_deq_bits_data(rob_io_deq_bits_data),
    .io_deq_bits_id(rob_io_deq_bits_id),
    .io_deq_bits_brAddr(rob_io_deq_bits_brAddr),
    .io_deq_bits_brTaken(rob_io_deq_bits_brTaken),
    .io_deq_bits_excpAddr(rob_io_deq_bits_excpAddr),
    .io_deq_bits_excpValid(rob_io_deq_bits_excpValid),
    .io_deq_bits_pc(rob_io_deq_bits_pc),
    .io_deq_bits_inst(rob_io_deq_bits_inst),
    .io_rs_0_valid(rob_io_rs_0_valid),
    .io_rs_0_bits_id(rob_io_rs_0_bits_id),
    .io_rs_1_valid(rob_io_rs_1_valid),
    .io_rs_1_bits_id(rob_io_rs_1_bits_id),
    .io_rs_2_valid(rob_io_rs_2_valid),
    .io_rs_2_bits_id(rob_io_rs_2_bits_id),
    .io_rs_3_valid(rob_io_rs_3_valid),
    .io_rs_3_bits_id(rob_io_rs_3_bits_id),
    .io_read_0_busy(rob_io_read_0_busy),
    .io_read_0_state(rob_io_read_0_state),
    .io_read_0_rd(rob_io_read_0_rd),
    .io_read_0_data(rob_io_read_0_data),
    .io_read_1_busy(rob_io_read_1_busy),
    .io_read_1_state(rob_io_read_1_state),
    .io_read_1_rd(rob_io_read_1_rd),
    .io_read_1_data(rob_io_read_1_data),
    .io_read_2_busy(rob_io_read_2_busy),
    .io_read_2_state(rob_io_read_2_state),
    .io_read_2_rd(rob_io_read_2_rd),
    .io_read_2_data(rob_io_read_2_data),
    .io_read_3_busy(rob_io_read_3_busy),
    .io_read_3_state(rob_io_read_3_state),
    .io_read_3_rd(rob_io_read_3_rd),
    .io_read_3_data(rob_io_read_3_data),
    .io_read_4_busy(rob_io_read_4_busy),
    .io_read_4_state(rob_io_read_4_state),
    .io_read_4_rd(rob_io_read_4_rd),
    .io_read_4_data(rob_io_read_4_data),
    .io_fu_0_valid(rob_io_fu_0_valid),
    .io_fu_0_bits_id(rob_io_fu_0_bits_id),
    .io_fu_0_bits_data(rob_io_fu_0_bits_data),
    .io_fu_1_valid(rob_io_fu_1_valid),
    .io_fu_1_bits_id(rob_io_fu_1_bits_id),
    .io_fu_1_bits_data(rob_io_fu_1_bits_data),
    .io_fu_1_bits_brAddr(rob_io_fu_1_bits_brAddr),
    .io_fu_1_bits_brTaken(rob_io_fu_1_bits_brTaken),
    .io_fu_2_valid(rob_io_fu_2_valid),
    .io_fu_2_bits_id(rob_io_fu_2_bits_id),
    .io_fu_2_bits_data(rob_io_fu_2_bits_data),
    .io_fu_3_valid(rob_io_fu_3_valid),
    .io_fu_3_bits_id(rob_io_fu_3_bits_id),
    .io_fu_3_bits_data(rob_io_fu_3_bits_data),
    .io_fu_3_bits_excpAddr(rob_io_fu_3_bits_excpAddr),
    .io_fu_3_bits_excpValid(rob_io_fu_3_bits_excpValid),
    .io_id(rob_io_id),
    .io_regStatus_0_owner(rob_io_regStatus_0_owner),
    .io_regStatus_1_owner(rob_io_regStatus_1_owner),
    .io_regStatus_2_owner(rob_io_regStatus_2_owner),
    .io_regStatus_3_owner(rob_io_regStatus_3_owner),
    .io_regStatus_4_owner(rob_io_regStatus_4_owner),
    .io_regStatus_5_owner(rob_io_regStatus_5_owner),
    .io_regStatus_6_owner(rob_io_regStatus_6_owner),
    .io_regStatus_7_owner(rob_io_regStatus_7_owner),
    .io_regStatus_8_owner(rob_io_regStatus_8_owner),
    .io_regStatus_9_owner(rob_io_regStatus_9_owner),
    .io_regStatus_10_owner(rob_io_regStatus_10_owner),
    .io_regStatus_11_owner(rob_io_regStatus_11_owner),
    .io_regStatus_12_owner(rob_io_regStatus_12_owner),
    .io_regStatus_13_owner(rob_io_regStatus_13_owner),
    .io_regStatus_14_owner(rob_io_regStatus_14_owner),
    .io_regStatus_15_owner(rob_io_regStatus_15_owner),
    .io_regStatus_16_owner(rob_io_regStatus_16_owner),
    .io_regStatus_17_owner(rob_io_regStatus_17_owner),
    .io_regStatus_18_owner(rob_io_regStatus_18_owner),
    .io_regStatus_19_owner(rob_io_regStatus_19_owner),
    .io_regStatus_20_owner(rob_io_regStatus_20_owner),
    .io_regStatus_21_owner(rob_io_regStatus_21_owner),
    .io_regStatus_22_owner(rob_io_regStatus_22_owner),
    .io_regStatus_23_owner(rob_io_regStatus_23_owner),
    .io_regStatus_24_owner(rob_io_regStatus_24_owner),
    .io_regStatus_25_owner(rob_io_regStatus_25_owner),
    .io_regStatus_26_owner(rob_io_regStatus_26_owner),
    .io_regStatus_27_owner(rob_io_regStatus_27_owner),
    .io_regStatus_28_owner(rob_io_regStatus_28_owner),
    .io_regStatus_29_owner(rob_io_regStatus_29_owner),
    .io_regStatus_30_owner(rob_io_regStatus_30_owner),
    .io_regStatus_31_owner(rob_io_regStatus_31_owner),
    .io_flush(rob_io_flush)
  );
  ALUStage_1 aluStage_1 ( // @[Core_1.scala 81:28]
    .clock(aluStage_1_clock),
    .reset(aluStage_1_reset),
    .io_in_ready(aluStage_1_io_in_ready),
    .io_in_valid(aluStage_1_io_in_valid),
    .io_in_bits_opr1(aluStage_1_io_in_bits_opr1),
    .io_in_bits_opr2(aluStage_1_io_in_bits_opr2),
    .io_in_bits_aluOp(aluStage_1_io_in_bits_aluOp),
    .io_in_bits_immSrc(aluStage_1_io_in_bits_immSrc),
    .io_in_bits_immSign(aluStage_1_io_in_bits_immSign),
    .io_in_bits_rs1Val(aluStage_1_io_in_bits_rs1Val),
    .io_in_bits_rs2Val(aluStage_1_io_in_bits_rs2Val),
    .io_in_bits_inst(aluStage_1_io_in_bits_inst),
    .io_in_bits_pc(aluStage_1_io_in_bits_pc),
    .io_in_bits_id(aluStage_1_io_in_bits_id),
    .io_out_valid(aluStage_1_io_out_valid),
    .io_out_bits_data(aluStage_1_io_out_bits_data),
    .io_out_bits_id(aluStage_1_io_out_bits_id),
    .io_out_bits_rd(aluStage_1_io_out_bits_rd),
    .io_flush(aluStage_1_io_flush)
  );
  ReservationStation aluRS ( // @[Core_1.scala 82:23]
    .clock(aluRS_clock),
    .reset(aluRS_reset),
    .io_enq_ready(aluRS_io_enq_ready),
    .io_enq_valid(aluRS_io_enq_valid),
    .io_enq_bits_op(aluRS_io_enq_bits_op),
    .io_enq_bits_opr1(aluRS_io_enq_bits_opr1),
    .io_enq_bits_opr2(aluRS_io_enq_bits_opr2),
    .io_enq_bits_rs1(aluRS_io_enq_bits_rs1),
    .io_enq_bits_rs2(aluRS_io_enq_bits_rs2),
    .io_enq_bits_ROBId(aluRS_io_enq_bits_ROBId),
    .io_enq_bits_rs1ROBId(aluRS_io_enq_bits_rs1ROBId),
    .io_enq_bits_rs2ROBId(aluRS_io_enq_bits_rs2ROBId),
    .io_enq_bits_immSrc(aluRS_io_enq_bits_immSrc),
    .io_enq_bits_immSign(aluRS_io_enq_bits_immSign),
    .io_enq_bits_excpType(aluRS_io_enq_bits_excpType),
    .io_enq_bits_pc(aluRS_io_enq_bits_pc),
    .io_enq_bits_inst(aluRS_io_enq_bits_inst),
    .io_deq_ready(aluRS_io_deq_ready),
    .io_deq_valid(aluRS_io_deq_valid),
    .io_deq_bits_op(aluRS_io_deq_bits_op),
    .io_deq_bits_ROBId(aluRS_io_deq_bits_ROBId),
    .io_deq_bits_opr1(aluRS_io_deq_bits_opr1),
    .io_deq_bits_opr2(aluRS_io_deq_bits_opr2),
    .io_deq_bits_rs1Val(aluRS_io_deq_bits_rs1Val),
    .io_deq_bits_rs2Val(aluRS_io_deq_bits_rs2Val),
    .io_deq_bits_immSrc(aluRS_io_deq_bits_immSrc),
    .io_deq_bits_immSign(aluRS_io_deq_bits_immSign),
    .io_deq_bits_excpType(aluRS_io_deq_bits_excpType),
    .io_deq_bits_pc(aluRS_io_deq_bits_pc),
    .io_deq_bits_inst(aluRS_io_deq_bits_inst),
    .io_robOut_valid(aluRS_io_robOut_valid),
    .io_robOut_bits_id(aluRS_io_robOut_bits_id),
    .io_robRead_0_busy(aluRS_io_robRead_0_busy),
    .io_robRead_0_state(aluRS_io_robRead_0_state),
    .io_robRead_0_rd(aluRS_io_robRead_0_rd),
    .io_robRead_0_data(aluRS_io_robRead_0_data),
    .io_robRead_1_busy(aluRS_io_robRead_1_busy),
    .io_robRead_1_state(aluRS_io_robRead_1_state),
    .io_robRead_1_rd(aluRS_io_robRead_1_rd),
    .io_robRead_1_data(aluRS_io_robRead_1_data),
    .io_robRead_2_busy(aluRS_io_robRead_2_busy),
    .io_robRead_2_state(aluRS_io_robRead_2_state),
    .io_robRead_2_rd(aluRS_io_robRead_2_rd),
    .io_robRead_2_data(aluRS_io_robRead_2_data),
    .io_robRead_3_busy(aluRS_io_robRead_3_busy),
    .io_robRead_3_state(aluRS_io_robRead_3_state),
    .io_robRead_3_rd(aluRS_io_robRead_3_rd),
    .io_robRead_3_data(aluRS_io_robRead_3_data),
    .io_robRead_4_busy(aluRS_io_robRead_4_busy),
    .io_robRead_4_state(aluRS_io_robRead_4_state),
    .io_robRead_4_rd(aluRS_io_robRead_4_rd),
    .io_robRead_4_data(aluRS_io_robRead_4_data),
    .io_regStatus_0_owner(aluRS_io_regStatus_0_owner),
    .io_regStatus_1_owner(aluRS_io_regStatus_1_owner),
    .io_regStatus_2_owner(aluRS_io_regStatus_2_owner),
    .io_regStatus_3_owner(aluRS_io_regStatus_3_owner),
    .io_regStatus_4_owner(aluRS_io_regStatus_4_owner),
    .io_regStatus_5_owner(aluRS_io_regStatus_5_owner),
    .io_regStatus_6_owner(aluRS_io_regStatus_6_owner),
    .io_regStatus_7_owner(aluRS_io_regStatus_7_owner),
    .io_regStatus_8_owner(aluRS_io_regStatus_8_owner),
    .io_regStatus_9_owner(aluRS_io_regStatus_9_owner),
    .io_regStatus_10_owner(aluRS_io_regStatus_10_owner),
    .io_regStatus_11_owner(aluRS_io_regStatus_11_owner),
    .io_regStatus_12_owner(aluRS_io_regStatus_12_owner),
    .io_regStatus_13_owner(aluRS_io_regStatus_13_owner),
    .io_regStatus_14_owner(aluRS_io_regStatus_14_owner),
    .io_regStatus_15_owner(aluRS_io_regStatus_15_owner),
    .io_regStatus_16_owner(aluRS_io_regStatus_16_owner),
    .io_regStatus_17_owner(aluRS_io_regStatus_17_owner),
    .io_regStatus_18_owner(aluRS_io_regStatus_18_owner),
    .io_regStatus_19_owner(aluRS_io_regStatus_19_owner),
    .io_regStatus_20_owner(aluRS_io_regStatus_20_owner),
    .io_regStatus_21_owner(aluRS_io_regStatus_21_owner),
    .io_regStatus_22_owner(aluRS_io_regStatus_22_owner),
    .io_regStatus_23_owner(aluRS_io_regStatus_23_owner),
    .io_regStatus_24_owner(aluRS_io_regStatus_24_owner),
    .io_regStatus_25_owner(aluRS_io_regStatus_25_owner),
    .io_regStatus_26_owner(aluRS_io_regStatus_26_owner),
    .io_regStatus_27_owner(aluRS_io_regStatus_27_owner),
    .io_regStatus_28_owner(aluRS_io_regStatus_28_owner),
    .io_regStatus_29_owner(aluRS_io_regStatus_29_owner),
    .io_regStatus_30_owner(aluRS_io_regStatus_30_owner),
    .io_regStatus_31_owner(aluRS_io_regStatus_31_owner),
    .io_cdb_0_valid(aluRS_io_cdb_0_valid),
    .io_cdb_0_bits_data(aluRS_io_cdb_0_bits_data),
    .io_cdb_0_bits_id(aluRS_io_cdb_0_bits_id),
    .io_cdb_0_bits_rd(aluRS_io_cdb_0_bits_rd),
    .io_cdb_1_valid(aluRS_io_cdb_1_valid),
    .io_cdb_1_bits_data(aluRS_io_cdb_1_bits_data),
    .io_cdb_1_bits_id(aluRS_io_cdb_1_bits_id),
    .io_cdb_1_bits_rd(aluRS_io_cdb_1_bits_rd),
    .io_cdb_2_valid(aluRS_io_cdb_2_valid),
    .io_cdb_2_bits_data(aluRS_io_cdb_2_bits_data),
    .io_cdb_2_bits_id(aluRS_io_cdb_2_bits_id),
    .io_cdb_2_bits_rd(aluRS_io_cdb_2_bits_rd),
    .io_cdb_3_valid(aluRS_io_cdb_3_valid),
    .io_cdb_3_bits_data(aluRS_io_cdb_3_bits_data),
    .io_cdb_3_bits_id(aluRS_io_cdb_3_bits_id),
    .io_cdb_3_bits_rd(aluRS_io_cdb_3_bits_rd),
    .io_rf_0_addr(aluRS_io_rf_0_addr),
    .io_rf_0_data(aluRS_io_rf_0_data),
    .io_rf_1_addr(aluRS_io_rf_1_addr),
    .io_rf_1_data(aluRS_io_rf_1_data),
    .io_flush(aluRS_io_flush)
  );
  BRUStage_1 bruStage_1 ( // @[Core_1.scala 84:28]
    .clock(bruStage_1_clock),
    .reset(bruStage_1_reset),
    .io_in_ready(bruStage_1_io_in_ready),
    .io_in_valid(bruStage_1_io_in_valid),
    .io_in_bits_opr1(bruStage_1_io_in_bits_opr1),
    .io_in_bits_opr2(bruStage_1_io_in_bits_opr2),
    .io_in_bits_bruOp(bruStage_1_io_in_bits_bruOp),
    .io_in_bits_immSrc(bruStage_1_io_in_bits_immSrc),
    .io_in_bits_rs1Val(bruStage_1_io_in_bits_rs1Val),
    .io_in_bits_rs2Val(bruStage_1_io_in_bits_rs2Val),
    .io_in_bits_inst(bruStage_1_io_in_bits_inst),
    .io_in_bits_pc(bruStage_1_io_in_bits_pc),
    .io_in_bits_id(bruStage_1_io_in_bits_id),
    .io_out_valid(bruStage_1_io_out_valid),
    .io_out_bits_brTaken(bruStage_1_io_out_bits_brTaken),
    .io_out_bits_brAddr(bruStage_1_io_out_bits_brAddr),
    .io_out_bits_rd(bruStage_1_io_out_bits_rd),
    .io_out_bits_data(bruStage_1_io_out_bits_data),
    .io_out_bits_id(bruStage_1_io_out_bits_id),
    .io_flush(bruStage_1_io_flush)
  );
  ReservationStation bruRS ( // @[Core_1.scala 85:23]
    .clock(bruRS_clock),
    .reset(bruRS_reset),
    .io_enq_ready(bruRS_io_enq_ready),
    .io_enq_valid(bruRS_io_enq_valid),
    .io_enq_bits_op(bruRS_io_enq_bits_op),
    .io_enq_bits_opr1(bruRS_io_enq_bits_opr1),
    .io_enq_bits_opr2(bruRS_io_enq_bits_opr2),
    .io_enq_bits_rs1(bruRS_io_enq_bits_rs1),
    .io_enq_bits_rs2(bruRS_io_enq_bits_rs2),
    .io_enq_bits_ROBId(bruRS_io_enq_bits_ROBId),
    .io_enq_bits_rs1ROBId(bruRS_io_enq_bits_rs1ROBId),
    .io_enq_bits_rs2ROBId(bruRS_io_enq_bits_rs2ROBId),
    .io_enq_bits_immSrc(bruRS_io_enq_bits_immSrc),
    .io_enq_bits_immSign(bruRS_io_enq_bits_immSign),
    .io_enq_bits_excpType(bruRS_io_enq_bits_excpType),
    .io_enq_bits_pc(bruRS_io_enq_bits_pc),
    .io_enq_bits_inst(bruRS_io_enq_bits_inst),
    .io_deq_ready(bruRS_io_deq_ready),
    .io_deq_valid(bruRS_io_deq_valid),
    .io_deq_bits_op(bruRS_io_deq_bits_op),
    .io_deq_bits_ROBId(bruRS_io_deq_bits_ROBId),
    .io_deq_bits_opr1(bruRS_io_deq_bits_opr1),
    .io_deq_bits_opr2(bruRS_io_deq_bits_opr2),
    .io_deq_bits_rs1Val(bruRS_io_deq_bits_rs1Val),
    .io_deq_bits_rs2Val(bruRS_io_deq_bits_rs2Val),
    .io_deq_bits_immSrc(bruRS_io_deq_bits_immSrc),
    .io_deq_bits_immSign(bruRS_io_deq_bits_immSign),
    .io_deq_bits_excpType(bruRS_io_deq_bits_excpType),
    .io_deq_bits_pc(bruRS_io_deq_bits_pc),
    .io_deq_bits_inst(bruRS_io_deq_bits_inst),
    .io_robOut_valid(bruRS_io_robOut_valid),
    .io_robOut_bits_id(bruRS_io_robOut_bits_id),
    .io_robRead_0_busy(bruRS_io_robRead_0_busy),
    .io_robRead_0_state(bruRS_io_robRead_0_state),
    .io_robRead_0_rd(bruRS_io_robRead_0_rd),
    .io_robRead_0_data(bruRS_io_robRead_0_data),
    .io_robRead_1_busy(bruRS_io_robRead_1_busy),
    .io_robRead_1_state(bruRS_io_robRead_1_state),
    .io_robRead_1_rd(bruRS_io_robRead_1_rd),
    .io_robRead_1_data(bruRS_io_robRead_1_data),
    .io_robRead_2_busy(bruRS_io_robRead_2_busy),
    .io_robRead_2_state(bruRS_io_robRead_2_state),
    .io_robRead_2_rd(bruRS_io_robRead_2_rd),
    .io_robRead_2_data(bruRS_io_robRead_2_data),
    .io_robRead_3_busy(bruRS_io_robRead_3_busy),
    .io_robRead_3_state(bruRS_io_robRead_3_state),
    .io_robRead_3_rd(bruRS_io_robRead_3_rd),
    .io_robRead_3_data(bruRS_io_robRead_3_data),
    .io_robRead_4_busy(bruRS_io_robRead_4_busy),
    .io_robRead_4_state(bruRS_io_robRead_4_state),
    .io_robRead_4_rd(bruRS_io_robRead_4_rd),
    .io_robRead_4_data(bruRS_io_robRead_4_data),
    .io_regStatus_0_owner(bruRS_io_regStatus_0_owner),
    .io_regStatus_1_owner(bruRS_io_regStatus_1_owner),
    .io_regStatus_2_owner(bruRS_io_regStatus_2_owner),
    .io_regStatus_3_owner(bruRS_io_regStatus_3_owner),
    .io_regStatus_4_owner(bruRS_io_regStatus_4_owner),
    .io_regStatus_5_owner(bruRS_io_regStatus_5_owner),
    .io_regStatus_6_owner(bruRS_io_regStatus_6_owner),
    .io_regStatus_7_owner(bruRS_io_regStatus_7_owner),
    .io_regStatus_8_owner(bruRS_io_regStatus_8_owner),
    .io_regStatus_9_owner(bruRS_io_regStatus_9_owner),
    .io_regStatus_10_owner(bruRS_io_regStatus_10_owner),
    .io_regStatus_11_owner(bruRS_io_regStatus_11_owner),
    .io_regStatus_12_owner(bruRS_io_regStatus_12_owner),
    .io_regStatus_13_owner(bruRS_io_regStatus_13_owner),
    .io_regStatus_14_owner(bruRS_io_regStatus_14_owner),
    .io_regStatus_15_owner(bruRS_io_regStatus_15_owner),
    .io_regStatus_16_owner(bruRS_io_regStatus_16_owner),
    .io_regStatus_17_owner(bruRS_io_regStatus_17_owner),
    .io_regStatus_18_owner(bruRS_io_regStatus_18_owner),
    .io_regStatus_19_owner(bruRS_io_regStatus_19_owner),
    .io_regStatus_20_owner(bruRS_io_regStatus_20_owner),
    .io_regStatus_21_owner(bruRS_io_regStatus_21_owner),
    .io_regStatus_22_owner(bruRS_io_regStatus_22_owner),
    .io_regStatus_23_owner(bruRS_io_regStatus_23_owner),
    .io_regStatus_24_owner(bruRS_io_regStatus_24_owner),
    .io_regStatus_25_owner(bruRS_io_regStatus_25_owner),
    .io_regStatus_26_owner(bruRS_io_regStatus_26_owner),
    .io_regStatus_27_owner(bruRS_io_regStatus_27_owner),
    .io_regStatus_28_owner(bruRS_io_regStatus_28_owner),
    .io_regStatus_29_owner(bruRS_io_regStatus_29_owner),
    .io_regStatus_30_owner(bruRS_io_regStatus_30_owner),
    .io_regStatus_31_owner(bruRS_io_regStatus_31_owner),
    .io_cdb_0_valid(bruRS_io_cdb_0_valid),
    .io_cdb_0_bits_data(bruRS_io_cdb_0_bits_data),
    .io_cdb_0_bits_id(bruRS_io_cdb_0_bits_id),
    .io_cdb_0_bits_rd(bruRS_io_cdb_0_bits_rd),
    .io_cdb_1_valid(bruRS_io_cdb_1_valid),
    .io_cdb_1_bits_data(bruRS_io_cdb_1_bits_data),
    .io_cdb_1_bits_id(bruRS_io_cdb_1_bits_id),
    .io_cdb_1_bits_rd(bruRS_io_cdb_1_bits_rd),
    .io_cdb_2_valid(bruRS_io_cdb_2_valid),
    .io_cdb_2_bits_data(bruRS_io_cdb_2_bits_data),
    .io_cdb_2_bits_id(bruRS_io_cdb_2_bits_id),
    .io_cdb_2_bits_rd(bruRS_io_cdb_2_bits_rd),
    .io_cdb_3_valid(bruRS_io_cdb_3_valid),
    .io_cdb_3_bits_data(bruRS_io_cdb_3_bits_data),
    .io_cdb_3_bits_id(bruRS_io_cdb_3_bits_id),
    .io_cdb_3_bits_rd(bruRS_io_cdb_3_bits_rd),
    .io_rf_0_addr(bruRS_io_rf_0_addr),
    .io_rf_0_data(bruRS_io_rf_0_data),
    .io_rf_1_addr(bruRS_io_rf_1_addr),
    .io_rf_1_data(bruRS_io_rf_1_data),
    .io_flush(bruRS_io_flush)
  );
  LSUStage_1 lsuStage_1 ( // @[Core_1.scala 87:28]
    .clock(lsuStage_1_clock),
    .reset(lsuStage_1_reset),
    .io_in_ready(lsuStage_1_io_in_ready),
    .io_in_valid(lsuStage_1_io_in_valid),
    .io_in_bits_lsuOp(lsuStage_1_io_in_bits_lsuOp),
    .io_in_bits_immSrc(lsuStage_1_io_in_bits_immSrc),
    .io_in_bits_rs1Val(lsuStage_1_io_in_bits_rs1Val),
    .io_in_bits_rs2Val(lsuStage_1_io_in_bits_rs2Val),
    .io_in_bits_inst(lsuStage_1_io_in_bits_inst),
    .io_in_bits_id(lsuStage_1_io_in_bits_id),
    .io_out_valid(lsuStage_1_io_out_valid),
    .io_out_bits_rd(lsuStage_1_io_out_bits_rd),
    .io_out_bits_data(lsuStage_1_io_out_bits_data),
    .io_out_bits_id(lsuStage_1_io_out_bits_id),
    .io_cache_read_req_ready(lsuStage_1_io_cache_read_req_ready),
    .io_cache_read_req_valid(lsuStage_1_io_cache_read_req_valid),
    .io_cache_read_req_bits_addr(lsuStage_1_io_cache_read_req_bits_addr),
    .io_cache_read_resp_ready(lsuStage_1_io_cache_read_resp_ready),
    .io_cache_read_resp_valid(lsuStage_1_io_cache_read_resp_valid),
    .io_cache_read_resp_bits_data(lsuStage_1_io_cache_read_resp_bits_data),
    .io_cache_write_req_ready(lsuStage_1_io_cache_write_req_ready),
    .io_cache_write_req_valid(lsuStage_1_io_cache_write_req_valid),
    .io_cache_write_req_bits_addr(lsuStage_1_io_cache_write_req_bits_addr),
    .io_cache_write_req_bits_data(lsuStage_1_io_cache_write_req_bits_data),
    .io_cache_write_req_bits_mask(lsuStage_1_io_cache_write_req_bits_mask),
    .io_cache_write_resp_ready(lsuStage_1_io_cache_write_resp_ready),
    .io_cache_write_resp_valid(lsuStage_1_io_cache_write_resp_valid),
    .io_rob_bits_id(lsuStage_1_io_rob_bits_id),
    .io_flush(lsuStage_1_io_flush)
  );
  ReservationStation lsuRS ( // @[Core_1.scala 88:23]
    .clock(lsuRS_clock),
    .reset(lsuRS_reset),
    .io_enq_ready(lsuRS_io_enq_ready),
    .io_enq_valid(lsuRS_io_enq_valid),
    .io_enq_bits_op(lsuRS_io_enq_bits_op),
    .io_enq_bits_opr1(lsuRS_io_enq_bits_opr1),
    .io_enq_bits_opr2(lsuRS_io_enq_bits_opr2),
    .io_enq_bits_rs1(lsuRS_io_enq_bits_rs1),
    .io_enq_bits_rs2(lsuRS_io_enq_bits_rs2),
    .io_enq_bits_ROBId(lsuRS_io_enq_bits_ROBId),
    .io_enq_bits_rs1ROBId(lsuRS_io_enq_bits_rs1ROBId),
    .io_enq_bits_rs2ROBId(lsuRS_io_enq_bits_rs2ROBId),
    .io_enq_bits_immSrc(lsuRS_io_enq_bits_immSrc),
    .io_enq_bits_immSign(lsuRS_io_enq_bits_immSign),
    .io_enq_bits_excpType(lsuRS_io_enq_bits_excpType),
    .io_enq_bits_pc(lsuRS_io_enq_bits_pc),
    .io_enq_bits_inst(lsuRS_io_enq_bits_inst),
    .io_deq_ready(lsuRS_io_deq_ready),
    .io_deq_valid(lsuRS_io_deq_valid),
    .io_deq_bits_op(lsuRS_io_deq_bits_op),
    .io_deq_bits_ROBId(lsuRS_io_deq_bits_ROBId),
    .io_deq_bits_opr1(lsuRS_io_deq_bits_opr1),
    .io_deq_bits_opr2(lsuRS_io_deq_bits_opr2),
    .io_deq_bits_rs1Val(lsuRS_io_deq_bits_rs1Val),
    .io_deq_bits_rs2Val(lsuRS_io_deq_bits_rs2Val),
    .io_deq_bits_immSrc(lsuRS_io_deq_bits_immSrc),
    .io_deq_bits_immSign(lsuRS_io_deq_bits_immSign),
    .io_deq_bits_excpType(lsuRS_io_deq_bits_excpType),
    .io_deq_bits_pc(lsuRS_io_deq_bits_pc),
    .io_deq_bits_inst(lsuRS_io_deq_bits_inst),
    .io_robOut_valid(lsuRS_io_robOut_valid),
    .io_robOut_bits_id(lsuRS_io_robOut_bits_id),
    .io_robRead_0_busy(lsuRS_io_robRead_0_busy),
    .io_robRead_0_state(lsuRS_io_robRead_0_state),
    .io_robRead_0_rd(lsuRS_io_robRead_0_rd),
    .io_robRead_0_data(lsuRS_io_robRead_0_data),
    .io_robRead_1_busy(lsuRS_io_robRead_1_busy),
    .io_robRead_1_state(lsuRS_io_robRead_1_state),
    .io_robRead_1_rd(lsuRS_io_robRead_1_rd),
    .io_robRead_1_data(lsuRS_io_robRead_1_data),
    .io_robRead_2_busy(lsuRS_io_robRead_2_busy),
    .io_robRead_2_state(lsuRS_io_robRead_2_state),
    .io_robRead_2_rd(lsuRS_io_robRead_2_rd),
    .io_robRead_2_data(lsuRS_io_robRead_2_data),
    .io_robRead_3_busy(lsuRS_io_robRead_3_busy),
    .io_robRead_3_state(lsuRS_io_robRead_3_state),
    .io_robRead_3_rd(lsuRS_io_robRead_3_rd),
    .io_robRead_3_data(lsuRS_io_robRead_3_data),
    .io_robRead_4_busy(lsuRS_io_robRead_4_busy),
    .io_robRead_4_state(lsuRS_io_robRead_4_state),
    .io_robRead_4_rd(lsuRS_io_robRead_4_rd),
    .io_robRead_4_data(lsuRS_io_robRead_4_data),
    .io_regStatus_0_owner(lsuRS_io_regStatus_0_owner),
    .io_regStatus_1_owner(lsuRS_io_regStatus_1_owner),
    .io_regStatus_2_owner(lsuRS_io_regStatus_2_owner),
    .io_regStatus_3_owner(lsuRS_io_regStatus_3_owner),
    .io_regStatus_4_owner(lsuRS_io_regStatus_4_owner),
    .io_regStatus_5_owner(lsuRS_io_regStatus_5_owner),
    .io_regStatus_6_owner(lsuRS_io_regStatus_6_owner),
    .io_regStatus_7_owner(lsuRS_io_regStatus_7_owner),
    .io_regStatus_8_owner(lsuRS_io_regStatus_8_owner),
    .io_regStatus_9_owner(lsuRS_io_regStatus_9_owner),
    .io_regStatus_10_owner(lsuRS_io_regStatus_10_owner),
    .io_regStatus_11_owner(lsuRS_io_regStatus_11_owner),
    .io_regStatus_12_owner(lsuRS_io_regStatus_12_owner),
    .io_regStatus_13_owner(lsuRS_io_regStatus_13_owner),
    .io_regStatus_14_owner(lsuRS_io_regStatus_14_owner),
    .io_regStatus_15_owner(lsuRS_io_regStatus_15_owner),
    .io_regStatus_16_owner(lsuRS_io_regStatus_16_owner),
    .io_regStatus_17_owner(lsuRS_io_regStatus_17_owner),
    .io_regStatus_18_owner(lsuRS_io_regStatus_18_owner),
    .io_regStatus_19_owner(lsuRS_io_regStatus_19_owner),
    .io_regStatus_20_owner(lsuRS_io_regStatus_20_owner),
    .io_regStatus_21_owner(lsuRS_io_regStatus_21_owner),
    .io_regStatus_22_owner(lsuRS_io_regStatus_22_owner),
    .io_regStatus_23_owner(lsuRS_io_regStatus_23_owner),
    .io_regStatus_24_owner(lsuRS_io_regStatus_24_owner),
    .io_regStatus_25_owner(lsuRS_io_regStatus_25_owner),
    .io_regStatus_26_owner(lsuRS_io_regStatus_26_owner),
    .io_regStatus_27_owner(lsuRS_io_regStatus_27_owner),
    .io_regStatus_28_owner(lsuRS_io_regStatus_28_owner),
    .io_regStatus_29_owner(lsuRS_io_regStatus_29_owner),
    .io_regStatus_30_owner(lsuRS_io_regStatus_30_owner),
    .io_regStatus_31_owner(lsuRS_io_regStatus_31_owner),
    .io_cdb_0_valid(lsuRS_io_cdb_0_valid),
    .io_cdb_0_bits_data(lsuRS_io_cdb_0_bits_data),
    .io_cdb_0_bits_id(lsuRS_io_cdb_0_bits_id),
    .io_cdb_0_bits_rd(lsuRS_io_cdb_0_bits_rd),
    .io_cdb_1_valid(lsuRS_io_cdb_1_valid),
    .io_cdb_1_bits_data(lsuRS_io_cdb_1_bits_data),
    .io_cdb_1_bits_id(lsuRS_io_cdb_1_bits_id),
    .io_cdb_1_bits_rd(lsuRS_io_cdb_1_bits_rd),
    .io_cdb_2_valid(lsuRS_io_cdb_2_valid),
    .io_cdb_2_bits_data(lsuRS_io_cdb_2_bits_data),
    .io_cdb_2_bits_id(lsuRS_io_cdb_2_bits_id),
    .io_cdb_2_bits_rd(lsuRS_io_cdb_2_bits_rd),
    .io_cdb_3_valid(lsuRS_io_cdb_3_valid),
    .io_cdb_3_bits_data(lsuRS_io_cdb_3_bits_data),
    .io_cdb_3_bits_id(lsuRS_io_cdb_3_bits_id),
    .io_cdb_3_bits_rd(lsuRS_io_cdb_3_bits_rd),
    .io_rf_0_addr(lsuRS_io_rf_0_addr),
    .io_rf_0_data(lsuRS_io_rf_0_data),
    .io_rf_1_addr(lsuRS_io_rf_1_addr),
    .io_rf_1_data(lsuRS_io_rf_1_data),
    .io_flush(lsuRS_io_flush)
  );
  CSRStage_1 csrStage_1 ( // @[Core_1.scala 90:28]
    .clock(csrStage_1_clock),
    .reset(csrStage_1_reset),
    .io_in_ready(csrStage_1_io_in_ready),
    .io_in_valid(csrStage_1_io_in_valid),
    .io_in_bits_csrOp(csrStage_1_io_in_bits_csrOp),
    .io_in_bits_excpType(csrStage_1_io_in_bits_excpType),
    .io_in_bits_rs1Val(csrStage_1_io_in_bits_rs1Val),
    .io_in_bits_inst(csrStage_1_io_in_bits_inst),
    .io_in_bits_id(csrStage_1_io_in_bits_id),
    .io_out_valid(csrStage_1_io_out_valid),
    .io_out_bits_rd(csrStage_1_io_out_bits_rd),
    .io_out_bits_data(csrStage_1_io_out_bits_data),
    .io_out_bits_excpAddr(csrStage_1_io_out_bits_excpAddr),
    .io_out_bits_excpValid(csrStage_1_io_out_bits_excpValid),
    .io_out_bits_id(csrStage_1_io_out_bits_id),
    .io_flush(csrStage_1_io_flush),
    .csrState_mcycle(csrStage_1_csrState_mcycle),
    .csrState_mcycleh(csrStage_1_csrState_mcycleh)
  );
  ReservationStation csrRS ( // @[Core_1.scala 91:23]
    .clock(csrRS_clock),
    .reset(csrRS_reset),
    .io_enq_ready(csrRS_io_enq_ready),
    .io_enq_valid(csrRS_io_enq_valid),
    .io_enq_bits_op(csrRS_io_enq_bits_op),
    .io_enq_bits_opr1(csrRS_io_enq_bits_opr1),
    .io_enq_bits_opr2(csrRS_io_enq_bits_opr2),
    .io_enq_bits_rs1(csrRS_io_enq_bits_rs1),
    .io_enq_bits_rs2(csrRS_io_enq_bits_rs2),
    .io_enq_bits_ROBId(csrRS_io_enq_bits_ROBId),
    .io_enq_bits_rs1ROBId(csrRS_io_enq_bits_rs1ROBId),
    .io_enq_bits_rs2ROBId(csrRS_io_enq_bits_rs2ROBId),
    .io_enq_bits_immSrc(csrRS_io_enq_bits_immSrc),
    .io_enq_bits_immSign(csrRS_io_enq_bits_immSign),
    .io_enq_bits_excpType(csrRS_io_enq_bits_excpType),
    .io_enq_bits_pc(csrRS_io_enq_bits_pc),
    .io_enq_bits_inst(csrRS_io_enq_bits_inst),
    .io_deq_ready(csrRS_io_deq_ready),
    .io_deq_valid(csrRS_io_deq_valid),
    .io_deq_bits_op(csrRS_io_deq_bits_op),
    .io_deq_bits_ROBId(csrRS_io_deq_bits_ROBId),
    .io_deq_bits_opr1(csrRS_io_deq_bits_opr1),
    .io_deq_bits_opr2(csrRS_io_deq_bits_opr2),
    .io_deq_bits_rs1Val(csrRS_io_deq_bits_rs1Val),
    .io_deq_bits_rs2Val(csrRS_io_deq_bits_rs2Val),
    .io_deq_bits_immSrc(csrRS_io_deq_bits_immSrc),
    .io_deq_bits_immSign(csrRS_io_deq_bits_immSign),
    .io_deq_bits_excpType(csrRS_io_deq_bits_excpType),
    .io_deq_bits_pc(csrRS_io_deq_bits_pc),
    .io_deq_bits_inst(csrRS_io_deq_bits_inst),
    .io_robOut_valid(csrRS_io_robOut_valid),
    .io_robOut_bits_id(csrRS_io_robOut_bits_id),
    .io_robRead_0_busy(csrRS_io_robRead_0_busy),
    .io_robRead_0_state(csrRS_io_robRead_0_state),
    .io_robRead_0_rd(csrRS_io_robRead_0_rd),
    .io_robRead_0_data(csrRS_io_robRead_0_data),
    .io_robRead_1_busy(csrRS_io_robRead_1_busy),
    .io_robRead_1_state(csrRS_io_robRead_1_state),
    .io_robRead_1_rd(csrRS_io_robRead_1_rd),
    .io_robRead_1_data(csrRS_io_robRead_1_data),
    .io_robRead_2_busy(csrRS_io_robRead_2_busy),
    .io_robRead_2_state(csrRS_io_robRead_2_state),
    .io_robRead_2_rd(csrRS_io_robRead_2_rd),
    .io_robRead_2_data(csrRS_io_robRead_2_data),
    .io_robRead_3_busy(csrRS_io_robRead_3_busy),
    .io_robRead_3_state(csrRS_io_robRead_3_state),
    .io_robRead_3_rd(csrRS_io_robRead_3_rd),
    .io_robRead_3_data(csrRS_io_robRead_3_data),
    .io_robRead_4_busy(csrRS_io_robRead_4_busy),
    .io_robRead_4_state(csrRS_io_robRead_4_state),
    .io_robRead_4_rd(csrRS_io_robRead_4_rd),
    .io_robRead_4_data(csrRS_io_robRead_4_data),
    .io_regStatus_0_owner(csrRS_io_regStatus_0_owner),
    .io_regStatus_1_owner(csrRS_io_regStatus_1_owner),
    .io_regStatus_2_owner(csrRS_io_regStatus_2_owner),
    .io_regStatus_3_owner(csrRS_io_regStatus_3_owner),
    .io_regStatus_4_owner(csrRS_io_regStatus_4_owner),
    .io_regStatus_5_owner(csrRS_io_regStatus_5_owner),
    .io_regStatus_6_owner(csrRS_io_regStatus_6_owner),
    .io_regStatus_7_owner(csrRS_io_regStatus_7_owner),
    .io_regStatus_8_owner(csrRS_io_regStatus_8_owner),
    .io_regStatus_9_owner(csrRS_io_regStatus_9_owner),
    .io_regStatus_10_owner(csrRS_io_regStatus_10_owner),
    .io_regStatus_11_owner(csrRS_io_regStatus_11_owner),
    .io_regStatus_12_owner(csrRS_io_regStatus_12_owner),
    .io_regStatus_13_owner(csrRS_io_regStatus_13_owner),
    .io_regStatus_14_owner(csrRS_io_regStatus_14_owner),
    .io_regStatus_15_owner(csrRS_io_regStatus_15_owner),
    .io_regStatus_16_owner(csrRS_io_regStatus_16_owner),
    .io_regStatus_17_owner(csrRS_io_regStatus_17_owner),
    .io_regStatus_18_owner(csrRS_io_regStatus_18_owner),
    .io_regStatus_19_owner(csrRS_io_regStatus_19_owner),
    .io_regStatus_20_owner(csrRS_io_regStatus_20_owner),
    .io_regStatus_21_owner(csrRS_io_regStatus_21_owner),
    .io_regStatus_22_owner(csrRS_io_regStatus_22_owner),
    .io_regStatus_23_owner(csrRS_io_regStatus_23_owner),
    .io_regStatus_24_owner(csrRS_io_regStatus_24_owner),
    .io_regStatus_25_owner(csrRS_io_regStatus_25_owner),
    .io_regStatus_26_owner(csrRS_io_regStatus_26_owner),
    .io_regStatus_27_owner(csrRS_io_regStatus_27_owner),
    .io_regStatus_28_owner(csrRS_io_regStatus_28_owner),
    .io_regStatus_29_owner(csrRS_io_regStatus_29_owner),
    .io_regStatus_30_owner(csrRS_io_regStatus_30_owner),
    .io_regStatus_31_owner(csrRS_io_regStatus_31_owner),
    .io_cdb_0_valid(csrRS_io_cdb_0_valid),
    .io_cdb_0_bits_data(csrRS_io_cdb_0_bits_data),
    .io_cdb_0_bits_id(csrRS_io_cdb_0_bits_id),
    .io_cdb_0_bits_rd(csrRS_io_cdb_0_bits_rd),
    .io_cdb_1_valid(csrRS_io_cdb_1_valid),
    .io_cdb_1_bits_data(csrRS_io_cdb_1_bits_data),
    .io_cdb_1_bits_id(csrRS_io_cdb_1_bits_id),
    .io_cdb_1_bits_rd(csrRS_io_cdb_1_bits_rd),
    .io_cdb_2_valid(csrRS_io_cdb_2_valid),
    .io_cdb_2_bits_data(csrRS_io_cdb_2_bits_data),
    .io_cdb_2_bits_id(csrRS_io_cdb_2_bits_id),
    .io_cdb_2_bits_rd(csrRS_io_cdb_2_bits_rd),
    .io_cdb_3_valid(csrRS_io_cdb_3_valid),
    .io_cdb_3_bits_data(csrRS_io_cdb_3_bits_data),
    .io_cdb_3_bits_id(csrRS_io_cdb_3_bits_id),
    .io_cdb_3_bits_rd(csrRS_io_cdb_3_bits_rd),
    .io_rf_0_addr(csrRS_io_rf_0_addr),
    .io_rf_0_data(csrRS_io_rf_0_data),
    .io_rf_1_addr(csrRS_io_rf_1_addr),
    .io_rf_1_data(csrRS_io_rf_1_data),
    .io_flush(csrRS_io_flush)
  );
  EdgeDetect edgeBackPressure ( // @[Core_1.scala 130:34]
    .clock(edgeBackPressure_clock),
    .io_in(edgeBackPressure_io_in),
    .io_change(edgeBackPressure_io_change)
  );
  Queue_5 fetch_pendingBranch ( // @[Core_1.scala 135:37]
    .clock(fetch_pendingBranch_clock),
    .reset(fetch_pendingBranch_reset),
    .io_enq_ready(fetch_pendingBranch_io_enq_ready),
    .io_enq_valid(fetch_pendingBranch_io_enq_valid),
    .io_enq_bits(fetch_pendingBranch_io_enq_bits),
    .io_deq_ready(fetch_pendingBranch_io_deq_ready),
    .io_deq_valid(fetch_pendingBranch_io_deq_valid),
    .io_deq_bits(fetch_pendingBranch_io_deq_bits)
  );
  Decoder_1 dec_decoders_0 ( // @[Core_1.scala 198:53]
    .io_inst(dec_decoders_0_io_inst),
    .io_out_brType(dec_decoders_0_io_out_brType),
    .io_out_wbType(dec_decoders_0_io_out_wbType),
    .io_out_lsuOp(dec_decoders_0_io_out_lsuOp),
    .io_out_aluOp(dec_decoders_0_io_out_aluOp),
    .io_out_opr1(dec_decoders_0_io_out_opr1),
    .io_out_opr2(dec_decoders_0_io_out_opr2),
    .io_out_immSrc(dec_decoders_0_io_out_immSrc),
    .io_out_immSign(dec_decoders_0_io_out_immSign),
    .io_out_csrOp(dec_decoders_0_io_out_csrOp),
    .io_out_excpType(dec_decoders_0_io_out_excpType)
  );
  Decoder_1 dec_decoders_1 ( // @[Core_1.scala 198:53]
    .io_inst(dec_decoders_1_io_inst),
    .io_out_brType(dec_decoders_1_io_out_brType),
    .io_out_wbType(dec_decoders_1_io_out_wbType),
    .io_out_lsuOp(dec_decoders_1_io_out_lsuOp),
    .io_out_aluOp(dec_decoders_1_io_out_aluOp),
    .io_out_opr1(dec_decoders_1_io_out_opr1),
    .io_out_opr2(dec_decoders_1_io_out_opr2),
    .io_out_immSrc(dec_decoders_1_io_out_immSrc),
    .io_out_immSign(dec_decoders_1_io_out_immSign),
    .io_out_csrOp(dec_decoders_1_io_out_csrOp),
    .io_out_excpType(dec_decoders_1_io_out_excpType)
  );
  Decoder_1 dec_decoders_2 ( // @[Core_1.scala 198:53]
    .io_inst(dec_decoders_2_io_inst),
    .io_out_brType(dec_decoders_2_io_out_brType),
    .io_out_wbType(dec_decoders_2_io_out_wbType),
    .io_out_lsuOp(dec_decoders_2_io_out_lsuOp),
    .io_out_aluOp(dec_decoders_2_io_out_aluOp),
    .io_out_opr1(dec_decoders_2_io_out_opr1),
    .io_out_opr2(dec_decoders_2_io_out_opr2),
    .io_out_immSrc(dec_decoders_2_io_out_immSrc),
    .io_out_immSign(dec_decoders_2_io_out_immSign),
    .io_out_csrOp(dec_decoders_2_io_out_csrOp),
    .io_out_excpType(dec_decoders_2_io_out_excpType)
  );
  Decoder_1 dec_decoders_3 ( // @[Core_1.scala 198:53]
    .io_inst(dec_decoders_3_io_inst),
    .io_out_brType(dec_decoders_3_io_out_brType),
    .io_out_wbType(dec_decoders_3_io_out_wbType),
    .io_out_lsuOp(dec_decoders_3_io_out_lsuOp),
    .io_out_aluOp(dec_decoders_3_io_out_aluOp),
    .io_out_opr1(dec_decoders_3_io_out_opr1),
    .io_out_opr2(dec_decoders_3_io_out_opr2),
    .io_out_immSrc(dec_decoders_3_io_out_immSrc),
    .io_out_immSign(dec_decoders_3_io_out_immSign),
    .io_out_csrOp(dec_decoders_3_io_out_csrOp),
    .io_out_excpType(dec_decoders_3_io_out_excpType)
  );
  DCache dcache ( // @[Core_1.scala 570:24]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_read_req_ready(dcache_io_read_req_ready),
    .io_read_req_valid(dcache_io_read_req_valid),
    .io_read_req_bits_addr(dcache_io_read_req_bits_addr),
    .io_read_resp_ready(dcache_io_read_resp_ready),
    .io_read_resp_valid(dcache_io_read_resp_valid),
    .io_read_resp_bits_data(dcache_io_read_resp_bits_data),
    .io_write_req_ready(dcache_io_write_req_ready),
    .io_write_req_valid(dcache_io_write_req_valid),
    .io_write_req_bits_addr(dcache_io_write_req_bits_addr),
    .io_write_req_bits_data(dcache_io_write_req_bits_data),
    .io_write_req_bits_mask(dcache_io_write_req_bits_mask),
    .io_write_resp_ready(dcache_io_write_resp_ready),
    .io_write_resp_valid(dcache_io_write_resp_valid),
    .io_tlbus_req_ready(dcache_io_tlbus_req_ready),
    .io_tlbus_req_valid(dcache_io_tlbus_req_valid),
    .io_tlbus_req_bits_opcode(dcache_io_tlbus_req_bits_opcode),
    .io_tlbus_req_bits_address(dcache_io_tlbus_req_bits_address),
    .io_tlbus_req_bits_data(dcache_io_tlbus_req_bits_data),
    .io_tlbus_resp_valid(dcache_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(dcache_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(dcache_io_tlbus_resp_bits_data),
    .io_flush(dcache_io_flush)
  );
  TLXbar xbar ( // @[Core_1.scala 695:22]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_masterFace_in_0_ready(xbar_io_masterFace_in_0_ready),
    .io_masterFace_in_0_valid(xbar_io_masterFace_in_0_valid),
    .io_masterFace_in_0_bits_address(xbar_io_masterFace_in_0_bits_address),
    .io_masterFace_in_1_ready(xbar_io_masterFace_in_1_ready),
    .io_masterFace_in_1_valid(xbar_io_masterFace_in_1_valid),
    .io_masterFace_in_1_bits_opcode(xbar_io_masterFace_in_1_bits_opcode),
    .io_masterFace_in_1_bits_address(xbar_io_masterFace_in_1_bits_address),
    .io_masterFace_in_1_bits_data(xbar_io_masterFace_in_1_bits_data),
    .io_masterFace_out_0_valid(xbar_io_masterFace_out_0_valid),
    .io_masterFace_out_0_bits_opcode(xbar_io_masterFace_out_0_bits_opcode),
    .io_masterFace_out_0_bits_data(xbar_io_masterFace_out_0_bits_data),
    .io_masterFace_out_1_valid(xbar_io_masterFace_out_1_valid),
    .io_masterFace_out_1_bits_opcode(xbar_io_masterFace_out_1_bits_opcode),
    .io_masterFace_out_1_bits_data(xbar_io_masterFace_out_1_bits_data),
    .io_slaveFace_in_0_ready(xbar_io_slaveFace_in_0_ready),
    .io_slaveFace_in_0_valid(xbar_io_slaveFace_in_0_valid),
    .io_slaveFace_in_0_bits_opcode(xbar_io_slaveFace_in_0_bits_opcode),
    .io_slaveFace_in_0_bits_size(xbar_io_slaveFace_in_0_bits_size),
    .io_slaveFace_in_0_bits_address(xbar_io_slaveFace_in_0_bits_address),
    .io_slaveFace_in_0_bits_data(xbar_io_slaveFace_in_0_bits_data),
    .io_slaveFace_out_0_ready(xbar_io_slaveFace_out_0_ready),
    .io_slaveFace_out_0_valid(xbar_io_slaveFace_out_0_valid),
    .io_slaveFace_out_0_bits_opcode(xbar_io_slaveFace_out_0_bits_opcode),
    .io_slaveFace_out_0_bits_data(xbar_io_slaveFace_out_0_bits_data)
  );
  SingleROM rom ( // @[Core_1.scala 696:21]
    .clock(rom_clock),
    .reset(rom_reset),
    .io_req_ready(rom_io_req_ready),
    .io_req_valid(rom_io_req_valid),
    .io_req_bits_opcode(rom_io_req_bits_opcode),
    .io_req_bits_size(rom_io_req_bits_size),
    .io_req_bits_address(rom_io_req_bits_address),
    .io_req_bits_data(rom_io_req_bits_data),
    .io_resp_ready(rom_io_resp_ready),
    .io_resp_valid(rom_io_resp_valid),
    .io_resp_bits_opcode(rom_io_resp_bits_opcode),
    .io_resp_bits_size(rom_io_resp_bits_size),
    .io_resp_bits_data(rom_io_resp_bits_data)
  );
  assign io_out_state_intRegState_regState_0 = rf_regState_0_regState_0; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_1 = rf_regState_0_regState_1; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_2 = rf_regState_0_regState_2; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_3 = rf_regState_0_regState_3; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_4 = rf_regState_0_regState_4; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_5 = rf_regState_0_regState_5; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_6 = rf_regState_0_regState_6; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_7 = rf_regState_0_regState_7; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_8 = rf_regState_0_regState_8; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_9 = rf_regState_0_regState_9; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_10 = rf_regState_0_regState_10; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_11 = rf_regState_0_regState_11; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_12 = rf_regState_0_regState_12; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_13 = rf_regState_0_regState_13; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_14 = rf_regState_0_regState_14; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_15 = rf_regState_0_regState_15; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_16 = rf_regState_0_regState_16; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_17 = rf_regState_0_regState_17; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_18 = rf_regState_0_regState_18; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_19 = rf_regState_0_regState_19; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_20 = rf_regState_0_regState_20; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_21 = rf_regState_0_regState_21; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_22 = rf_regState_0_regState_22; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_23 = rf_regState_0_regState_23; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_24 = rf_regState_0_regState_24; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_25 = rf_regState_0_regState_25; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_26 = rf_regState_0_regState_26; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_27 = rf_regState_0_regState_27; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_28 = rf_regState_0_regState_28; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_29 = rf_regState_0_regState_29; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_30 = rf_regState_0_regState_30; // @[Core_1.scala 681:28]
  assign io_out_state_intRegState_regState_31 = rf_regState_0_regState_31; // @[Core_1.scala 681:28]
  assign io_out_state_instState_commit = io_out_state_instState_REG_commit; // @[Core_1.scala 687:28]
  assign io_out_state_instState_pc = io_out_state_instState_REG_pc; // @[Core_1.scala 687:28]
  assign io_out_state_instState_inst = io_out_state_instState_REG_inst; // @[Core_1.scala 687:28]
  assign io_out_state_csrState_mcycle = csrStage_1_csrState_mcycle; // @[Core_1.scala 684:28]
  assign io_out_state_csrState_mcycleh = csrStage_1_csrState_mcycleh; // @[Core_1.scala 684:28]
  assign ib_clock = clock;
  assign ib_reset = reset;
  assign ib_io_in_valid = fetch_fire & (~blockValid | willWakeUp) & ~willBlock; // @[Core_1.scala 172:66]
  assign ib_io_in_bits_icache_data = icache_io_read_resp_bits_data; // @[Core_1.scala 173:26]
  assign ib_io_in_bits_icache_addr = icache_io_read_resp_bits_addr; // @[Core_1.scala 173:26]
  assign ib_io_in_bits_icache_inst_0 = icache_io_read_resp_bits_inst_0; // @[Core_1.scala 173:26]
  assign ib_io_in_bits_icache_inst_1 = icache_io_read_resp_bits_inst_1; // @[Core_1.scala 173:26]
  assign ib_io_in_bits_icache_inst_2 = icache_io_read_resp_bits_inst_2; // @[Core_1.scala 173:26]
  assign ib_io_in_bits_icache_inst_3 = icache_io_read_resp_bits_inst_3; // @[Core_1.scala 173:26]
  assign ib_io_in_bits_icache_size = icacheRespIsAlignAddr ? icache_io_read_resp_bits_size :
    _ib_io_in_bits_icache_size_T_2; // @[Core_1.scala 177:37]
  assign ib_io_in_bits_pc = icache_io_read_resp_bits_addr; // @[Core_1.scala 178:22]
  assign ib_io_in_bits_flush = globalBrTaken | reset; // @[Core_1.scala 179:42]
  assign ib_io_out_ready = ~dec_full | dec_fire; // @[Core_1.scala 193:28]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_read_req_valid = preFetchInst & io_in_start; // @[Core_1.scala 150:46]
  assign icache_io_read_req_bits_addr = _lastPc_T ? _icache_io_read_req_bits_addr_T_1 :
    _icache_io_read_req_bits_addr_T_2; // @[Core_1.scala 151:40]
  assign icache_io_read_resp_ready = ib_io_in_ready; // @[Core_1.scala 152:31]
  assign icache_io_tlbus_req_ready = xbar_io_masterFace_in_0_ready; // @[Core_1.scala 698:25]
  assign icache_io_tlbus_resp_valid = xbar_io_masterFace_out_0_valid; // @[Core_1.scala 699:26]
  assign icache_io_tlbus_resp_bits_opcode = xbar_io_masterFace_out_0_bits_opcode; // @[Core_1.scala 699:26]
  assign icache_io_tlbus_resp_bits_data = xbar_io_masterFace_out_0_bits_data; // @[Core_1.scala 699:26]
  assign icache_io_flush = globalBrTaken; // @[Core_1.scala 153:21]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_r_0_addr = aluRS_io_rf_0_addr; // @[Core_1.scala 651:20]
  assign rf_io_r_1_addr = aluRS_io_rf_1_addr; // @[Core_1.scala 652:20]
  assign rf_io_r_2_addr = bruRS_io_rf_0_addr; // @[Core_1.scala 653:20]
  assign rf_io_r_3_addr = bruRS_io_rf_1_addr; // @[Core_1.scala 654:20]
  assign rf_io_r_4_addr = lsuRS_io_rf_0_addr; // @[Core_1.scala 655:20]
  assign rf_io_r_5_addr = lsuRS_io_rf_1_addr; // @[Core_1.scala 656:20]
  assign rf_io_r_6_addr = csrRS_io_rf_0_addr; // @[Core_1.scala 657:20]
  assign rf_io_r_7_addr = csrRS_io_rf_1_addr; // @[Core_1.scala 658:20]
  assign rf_io_w_0_addr = rob_io_deq_bits_rd; // @[Core_1.scala 668:21]
  assign rf_io_w_0_en = rob_io_deq_bits_rdWrEn & _csrExcpValid_T; // @[Core_1.scala 670:45]
  assign rf_io_w_0_data = rob_io_deq_bits_data; // @[Core_1.scala 669:21]
  assign rob_clock = clock;
  assign rob_reset = reset;
  assign rob_io_enq_valid = (issue_aluValid | issue_bruValid | issue_lsuValid | issue_csrValid) & issue_full & rsReady; // @[Core_1.scala 462:110]
  assign rob_io_enq_bits_rd = invalidRd ? 5'h0 : rd; // @[Core_1.scala 477:23]
  assign rob_io_enq_bits_fuValid = {rob_io_enq_bits_fuValid_hi,rob_io_enq_bits_fuValid_lo}; // @[Cat.scala 33:92]
  assign rob_io_enq_bits_fuOp = {{3'd0}, _rob_io_enq_bits_fuOp_T_3}; // @[Core_1.scala 463:26]
  assign rob_io_enq_bits_pc = issue_stagePc; // @[Core_1.scala 471:24]
  assign rob_io_enq_bits_inst = _issue_chosenInst_T_10 | _issue_chosenInst_T_8; // @[Mux.scala 27:73]
  assign rob_io_deq_ready = 1'h1; // @[Core_1.scala 627:22]
  assign rob_io_rs_0_valid = aluRS_io_robOut_valid; // @[Core_1.scala 600:20]
  assign rob_io_rs_0_bits_id = aluRS_io_robOut_bits_id; // @[Core_1.scala 600:20]
  assign rob_io_rs_1_valid = bruRS_io_robOut_valid; // @[Core_1.scala 609:20]
  assign rob_io_rs_1_bits_id = bruRS_io_robOut_bits_id; // @[Core_1.scala 609:20]
  assign rob_io_rs_2_valid = lsuRS_io_robOut_valid; // @[Core_1.scala 616:20]
  assign rob_io_rs_2_bits_id = lsuRS_io_robOut_bits_id; // @[Core_1.scala 616:20]
  assign rob_io_rs_3_valid = csrRS_io_robOut_valid; // @[Core_1.scala 625:20]
  assign rob_io_rs_3_bits_id = csrRS_io_robOut_bits_id; // @[Core_1.scala 625:20]
  assign rob_io_fu_0_valid = aluStage_1_io_out_valid; // @[Core_1.scala 595:26]
  assign rob_io_fu_0_bits_id = aluStage_1_io_out_bits_id[2:0]; // @[Core_1.scala 598:28]
  assign rob_io_fu_0_bits_data = aluStage_1_io_out_bits_data; // @[Core_1.scala 597:30]
  assign rob_io_fu_1_valid = bruStage_1_io_out_valid; // @[Core_1.scala 602:26]
  assign rob_io_fu_1_bits_id = bruStage_1_io_out_bits_id[2:0]; // @[Core_1.scala 605:28]
  assign rob_io_fu_1_bits_data = bruStage_1_io_out_bits_data; // @[Core_1.scala 604:30]
  assign rob_io_fu_1_bits_brAddr = bruStage_1_io_out_bits_brAddr; // @[Core_1.scala 607:32]
  assign rob_io_fu_1_bits_brTaken = bruStage_1_io_out_bits_brTaken; // @[Core_1.scala 608:33]
  assign rob_io_fu_2_valid = lsuStage_1_io_out_valid; // @[Core_1.scala 611:26]
  assign rob_io_fu_2_bits_id = lsuStage_1_io_out_bits_id[2:0]; // @[Core_1.scala 614:28]
  assign rob_io_fu_2_bits_data = lsuStage_1_io_out_bits_data; // @[Core_1.scala 613:30]
  assign rob_io_fu_3_valid = csrStage_1_io_out_valid; // @[Core_1.scala 618:26]
  assign rob_io_fu_3_bits_id = csrStage_1_io_out_bits_id[2:0]; // @[Core_1.scala 621:28]
  assign rob_io_fu_3_bits_data = csrStage_1_io_out_bits_data; // @[Core_1.scala 620:30]
  assign rob_io_fu_3_bits_excpAddr = csrStage_1_io_out_bits_excpAddr; // @[Core_1.scala 624:34]
  assign rob_io_fu_3_bits_excpValid = csrStage_1_io_out_bits_excpValid; // @[Core_1.scala 623:35]
  assign rob_io_flush = globalBrTaken | reset; // @[Core_1.scala 479:35]
  assign aluStage_1_clock = clock;
  assign aluStage_1_reset = reset;
  assign aluStage_1_io_in_valid = aluRS_io_deq_valid; // @[Core_1.scala 511:28]
  assign aluStage_1_io_in_bits_opr1 = aluRS_io_deq_bits_opr1; // @[Core_1.scala 517:32]
  assign aluStage_1_io_in_bits_opr2 = aluRS_io_deq_bits_opr2; // @[Core_1.scala 518:32]
  assign aluStage_1_io_in_bits_aluOp = aluRS_io_deq_bits_op[4:0]; // @[Core_1.scala 512:33]
  assign aluStage_1_io_in_bits_immSrc = aluRS_io_deq_bits_immSrc; // @[Core_1.scala 513:34]
  assign aluStage_1_io_in_bits_immSign = aluRS_io_deq_bits_immSign; // @[Core_1.scala 514:35]
  assign aluStage_1_io_in_bits_rs1Val = aluRS_io_deq_bits_rs1Val; // @[Core_1.scala 520:34]
  assign aluStage_1_io_in_bits_rs2Val = aluRS_io_deq_bits_rs2Val; // @[Core_1.scala 521:34]
  assign aluStage_1_io_in_bits_inst = aluRS_io_deq_bits_inst; // @[Core_1.scala 515:32]
  assign aluStage_1_io_in_bits_pc = aluRS_io_deq_bits_pc; // @[Core_1.scala 516:30]
  assign aluStage_1_io_in_bits_id = aluRS_io_deq_bits_ROBId; // @[Core_1.scala 519:30]
  assign aluStage_1_io_flush = globalBrTaken | reset; // @[Core_1.scala 522:42]
  assign aluRS_clock = clock;
  assign aluRS_reset = reset;
  assign aluRS_io_enq_valid = issue_instFire & issue_aluValid; // @[Core_1.scala 505:43]
  assign aluRS_io_enq_bits_op = {{3'd0}, _rob_io_enq_bits_fuOp_T_3}; // @[Core_1.scala 482:23 489:16]
  assign aluRS_io_enq_bits_opr1 = _issue_chosenDecodesigs_T_45 | _issue_chosenDecodesigs_T_43; // @[Mux.scala 27:73]
  assign aluRS_io_enq_bits_opr2 = _issue_chosenDecodesigs_T_38 | _issue_chosenDecodesigs_T_36; // @[Mux.scala 27:73]
  assign aluRS_io_enq_bits_rs1 = issue_chosenDecodesigs_opr1 == 4'h1 ? rs1 : 5'h0; // @[Core_1.scala 266:24]
  assign aluRS_io_enq_bits_rs2 = issue_chosenDecodesigs_opr2 == 4'h2 ? rs2 : 5'h0; // @[Core_1.scala 267:24]
  assign aluRS_io_enq_bits_ROBId = {{5'd0}, rob_io_id}; // @[Core_1.scala 482:23 483:19]
  assign aluRS_io_enq_bits_rs1ROBId = 5'h1f == issue_rs1 ? rob_io_regStatus_31_owner : _GEN_106; // @[Core_1.scala 500:{22,22}]
  assign aluRS_io_enq_bits_rs2ROBId = 5'h1f == issue_rs1 ? rob_io_regStatus_31_owner : _GEN_106; // @[Core_1.scala 500:{22,22}]
  assign aluRS_io_enq_bits_immSrc = _issue_chosenDecodesigs_T_31 | _issue_chosenDecodesigs_T_29; // @[Mux.scala 27:73]
  assign aluRS_io_enq_bits_immSign = _issue_chosenDecodesigs_T[0] & issue_decodeSigs_0_immSign |
    _issue_chosenDecodesigs_T[1] & issue_decodeSigs_1_immSign | _issue_chosenDecodesigs_T[2] &
    issue_decodeSigs_2_immSign | _issue_chosenDecodesigs_T[3] & issue_decodeSigs_3_immSign; // @[Mux.scala 27:73]
  assign aluRS_io_enq_bits_excpType = _issue_chosenDecodesigs_T_10 | _issue_chosenDecodesigs_T_8; // @[Mux.scala 27:73]
  assign aluRS_io_enq_bits_pc = issue_stagePc; // @[Core_1.scala 482:23 488:16]
  assign aluRS_io_enq_bits_inst = _issue_chosenInst_T_10 | _issue_chosenInst_T_8; // @[Mux.scala 27:73]
  assign aluRS_io_deq_ready = aluStage_1_io_in_ready; // @[Core_1.scala 509:24]
  assign aluRS_io_robRead_0_busy = rob_io_read_0_busy; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_0_state = rob_io_read_0_state; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_0_rd = rob_io_read_0_rd; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_0_data = rob_io_read_0_data; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_1_busy = rob_io_read_1_busy; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_1_state = rob_io_read_1_state; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_1_rd = rob_io_read_1_rd; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_1_data = rob_io_read_1_data; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_2_busy = rob_io_read_2_busy; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_2_state = rob_io_read_2_state; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_2_rd = rob_io_read_2_rd; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_2_data = rob_io_read_2_data; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_3_busy = rob_io_read_3_busy; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_3_state = rob_io_read_3_state; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_3_rd = rob_io_read_3_rd; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_3_data = rob_io_read_3_data; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_4_busy = rob_io_read_4_busy; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_4_state = rob_io_read_4_state; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_4_rd = rob_io_read_4_rd; // @[Core_1.scala 646:16]
  assign aluRS_io_robRead_4_data = rob_io_read_4_data; // @[Core_1.scala 646:16]
  assign aluRS_io_regStatus_0_owner = rob_io_regStatus_0_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_1_owner = rob_io_regStatus_1_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_2_owner = rob_io_regStatus_2_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_3_owner = rob_io_regStatus_3_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_4_owner = rob_io_regStatus_4_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_5_owner = rob_io_regStatus_5_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_6_owner = rob_io_regStatus_6_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_7_owner = rob_io_regStatus_7_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_8_owner = rob_io_regStatus_8_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_9_owner = rob_io_regStatus_9_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_10_owner = rob_io_regStatus_10_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_11_owner = rob_io_regStatus_11_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_12_owner = rob_io_regStatus_12_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_13_owner = rob_io_regStatus_13_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_14_owner = rob_io_regStatus_14_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_15_owner = rob_io_regStatus_15_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_16_owner = rob_io_regStatus_16_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_17_owner = rob_io_regStatus_17_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_18_owner = rob_io_regStatus_18_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_19_owner = rob_io_regStatus_19_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_20_owner = rob_io_regStatus_20_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_21_owner = rob_io_regStatus_21_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_22_owner = rob_io_regStatus_22_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_23_owner = rob_io_regStatus_23_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_24_owner = rob_io_regStatus_24_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_25_owner = rob_io_regStatus_25_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_26_owner = rob_io_regStatus_26_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_27_owner = rob_io_regStatus_27_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_28_owner = rob_io_regStatus_28_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_29_owner = rob_io_regStatus_29_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_30_owner = rob_io_regStatus_30_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_regStatus_31_owner = rob_io_regStatus_31_owner; // @[Core_1.scala 507:24]
  assign aluRS_io_cdb_0_valid = aluStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign aluRS_io_cdb_0_bits_data = aluStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign aluRS_io_cdb_0_bits_id = aluStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign aluRS_io_cdb_0_bits_rd = aluStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign aluRS_io_cdb_1_valid = bruStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign aluRS_io_cdb_1_bits_data = bruStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign aluRS_io_cdb_1_bits_id = bruStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign aluRS_io_cdb_1_bits_rd = bruStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign aluRS_io_cdb_2_valid = lsuStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign aluRS_io_cdb_2_bits_data = lsuStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign aluRS_io_cdb_2_bits_id = lsuStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign aluRS_io_cdb_2_bits_rd = lsuStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign aluRS_io_cdb_3_valid = csrStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign aluRS_io_cdb_3_bits_data = csrStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign aluRS_io_cdb_3_bits_id = csrStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign aluRS_io_cdb_3_bits_rd = csrStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign aluRS_io_rf_0_data = rf_io_r_0_data; // @[Core_1.scala 651:20]
  assign aluRS_io_rf_1_data = rf_io_r_1_data; // @[Core_1.scala 652:20]
  assign aluRS_io_flush = globalBrTaken | reset; // @[Core_1.scala 508:37]
  assign bruStage_1_clock = clock;
  assign bruStage_1_reset = reset;
  assign bruStage_1_io_in_valid = bruRS_io_deq_valid; // @[Core_1.scala 534:28]
  assign bruStage_1_io_in_bits_opr1 = bruRS_io_deq_bits_opr1; // @[Core_1.scala 539:32]
  assign bruStage_1_io_in_bits_opr2 = bruRS_io_deq_bits_opr2; // @[Core_1.scala 540:32]
  assign bruStage_1_io_in_bits_bruOp = bruRS_io_deq_bits_op[3:0]; // @[Core_1.scala 535:33]
  assign bruStage_1_io_in_bits_immSrc = bruRS_io_deq_bits_immSrc; // @[Core_1.scala 536:34]
  assign bruStage_1_io_in_bits_rs1Val = bruRS_io_deq_bits_rs1Val; // @[Core_1.scala 542:34]
  assign bruStage_1_io_in_bits_rs2Val = bruRS_io_deq_bits_rs2Val; // @[Core_1.scala 543:34]
  assign bruStage_1_io_in_bits_inst = bruRS_io_deq_bits_inst; // @[Core_1.scala 537:32]
  assign bruStage_1_io_in_bits_pc = bruRS_io_deq_bits_pc; // @[Core_1.scala 538:30]
  assign bruStage_1_io_in_bits_id = bruRS_io_deq_bits_ROBId; // @[Core_1.scala 541:30]
  assign bruStage_1_io_flush = globalBrTaken | reset; // @[Core_1.scala 544:42]
  assign bruRS_clock = clock;
  assign bruRS_reset = reset;
  assign bruRS_io_enq_valid = issue_instFire & issue_bruValid; // @[Core_1.scala 528:43]
  assign bruRS_io_enq_bits_op = {{3'd0}, _rob_io_enq_bits_fuOp_T_3}; // @[Core_1.scala 482:23 489:16]
  assign bruRS_io_enq_bits_opr1 = _issue_chosenDecodesigs_T_45 | _issue_chosenDecodesigs_T_43; // @[Mux.scala 27:73]
  assign bruRS_io_enq_bits_opr2 = _issue_chosenDecodesigs_T_38 | _issue_chosenDecodesigs_T_36; // @[Mux.scala 27:73]
  assign bruRS_io_enq_bits_rs1 = issue_chosenDecodesigs_opr1 == 4'h1 ? rs1 : 5'h0; // @[Core_1.scala 266:24]
  assign bruRS_io_enq_bits_rs2 = issue_chosenDecodesigs_opr2 == 4'h2 ? rs2 : 5'h0; // @[Core_1.scala 267:24]
  assign bruRS_io_enq_bits_ROBId = {{5'd0}, rob_io_id}; // @[Core_1.scala 482:23 483:19]
  assign bruRS_io_enq_bits_rs1ROBId = 5'h1f == issue_rs1 ? rob_io_regStatus_31_owner : _GEN_106; // @[Core_1.scala 500:{22,22}]
  assign bruRS_io_enq_bits_rs2ROBId = 5'h1f == issue_rs1 ? rob_io_regStatus_31_owner : _GEN_106; // @[Core_1.scala 500:{22,22}]
  assign bruRS_io_enq_bits_immSrc = _issue_chosenDecodesigs_T_31 | _issue_chosenDecodesigs_T_29; // @[Mux.scala 27:73]
  assign bruRS_io_enq_bits_immSign = _issue_chosenDecodesigs_T[0] & issue_decodeSigs_0_immSign |
    _issue_chosenDecodesigs_T[1] & issue_decodeSigs_1_immSign | _issue_chosenDecodesigs_T[2] &
    issue_decodeSigs_2_immSign | _issue_chosenDecodesigs_T[3] & issue_decodeSigs_3_immSign; // @[Mux.scala 27:73]
  assign bruRS_io_enq_bits_excpType = _issue_chosenDecodesigs_T_10 | _issue_chosenDecodesigs_T_8; // @[Mux.scala 27:73]
  assign bruRS_io_enq_bits_pc = issue_stagePc; // @[Core_1.scala 482:23 488:16]
  assign bruRS_io_enq_bits_inst = _issue_chosenInst_T_10 | _issue_chosenInst_T_8; // @[Mux.scala 27:73]
  assign bruRS_io_deq_ready = bruStage_1_io_in_ready; // @[Core_1.scala 532:24]
  assign bruRS_io_robRead_0_busy = rob_io_read_0_busy; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_0_state = rob_io_read_0_state; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_0_rd = rob_io_read_0_rd; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_0_data = rob_io_read_0_data; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_1_busy = rob_io_read_1_busy; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_1_state = rob_io_read_1_state; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_1_rd = rob_io_read_1_rd; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_1_data = rob_io_read_1_data; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_2_busy = rob_io_read_2_busy; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_2_state = rob_io_read_2_state; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_2_rd = rob_io_read_2_rd; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_2_data = rob_io_read_2_data; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_3_busy = rob_io_read_3_busy; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_3_state = rob_io_read_3_state; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_3_rd = rob_io_read_3_rd; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_3_data = rob_io_read_3_data; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_4_busy = rob_io_read_4_busy; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_4_state = rob_io_read_4_state; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_4_rd = rob_io_read_4_rd; // @[Core_1.scala 646:16]
  assign bruRS_io_robRead_4_data = rob_io_read_4_data; // @[Core_1.scala 646:16]
  assign bruRS_io_regStatus_0_owner = rob_io_regStatus_0_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_1_owner = rob_io_regStatus_1_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_2_owner = rob_io_regStatus_2_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_3_owner = rob_io_regStatus_3_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_4_owner = rob_io_regStatus_4_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_5_owner = rob_io_regStatus_5_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_6_owner = rob_io_regStatus_6_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_7_owner = rob_io_regStatus_7_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_8_owner = rob_io_regStatus_8_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_9_owner = rob_io_regStatus_9_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_10_owner = rob_io_regStatus_10_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_11_owner = rob_io_regStatus_11_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_12_owner = rob_io_regStatus_12_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_13_owner = rob_io_regStatus_13_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_14_owner = rob_io_regStatus_14_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_15_owner = rob_io_regStatus_15_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_16_owner = rob_io_regStatus_16_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_17_owner = rob_io_regStatus_17_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_18_owner = rob_io_regStatus_18_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_19_owner = rob_io_regStatus_19_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_20_owner = rob_io_regStatus_20_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_21_owner = rob_io_regStatus_21_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_22_owner = rob_io_regStatus_22_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_23_owner = rob_io_regStatus_23_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_24_owner = rob_io_regStatus_24_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_25_owner = rob_io_regStatus_25_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_26_owner = rob_io_regStatus_26_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_27_owner = rob_io_regStatus_27_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_28_owner = rob_io_regStatus_28_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_29_owner = rob_io_regStatus_29_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_30_owner = rob_io_regStatus_30_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_regStatus_31_owner = rob_io_regStatus_31_owner; // @[Core_1.scala 530:24]
  assign bruRS_io_cdb_0_valid = aluStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign bruRS_io_cdb_0_bits_data = aluStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign bruRS_io_cdb_0_bits_id = aluStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign bruRS_io_cdb_0_bits_rd = aluStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign bruRS_io_cdb_1_valid = bruStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign bruRS_io_cdb_1_bits_data = bruStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign bruRS_io_cdb_1_bits_id = bruStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign bruRS_io_cdb_1_bits_rd = bruStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign bruRS_io_cdb_2_valid = lsuStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign bruRS_io_cdb_2_bits_data = lsuStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign bruRS_io_cdb_2_bits_id = lsuStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign bruRS_io_cdb_2_bits_rd = lsuStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign bruRS_io_cdb_3_valid = csrStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign bruRS_io_cdb_3_bits_data = csrStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign bruRS_io_cdb_3_bits_id = csrStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign bruRS_io_cdb_3_bits_rd = csrStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign bruRS_io_rf_0_data = rf_io_r_2_data; // @[Core_1.scala 653:20]
  assign bruRS_io_rf_1_data = rf_io_r_3_data; // @[Core_1.scala 654:20]
  assign bruRS_io_flush = globalBrTaken | reset; // @[Core_1.scala 531:37]
  assign lsuStage_1_clock = clock;
  assign lsuStage_1_reset = reset;
  assign lsuStage_1_io_in_valid = lsuRS_io_deq_valid; // @[Core_1.scala 555:28]
  assign lsuStage_1_io_in_bits_lsuOp = lsuRS_io_deq_bits_op[4:0]; // @[Core_1.scala 556:33]
  assign lsuStage_1_io_in_bits_immSrc = lsuRS_io_deq_bits_immSrc; // @[Core_1.scala 557:34]
  assign lsuStage_1_io_in_bits_rs1Val = lsuRS_io_deq_bits_rs1Val; // @[Core_1.scala 560:34]
  assign lsuStage_1_io_in_bits_rs2Val = lsuRS_io_deq_bits_rs2Val; // @[Core_1.scala 561:34]
  assign lsuStage_1_io_in_bits_inst = lsuRS_io_deq_bits_inst; // @[Core_1.scala 558:32]
  assign lsuStage_1_io_in_bits_id = lsuRS_io_deq_bits_ROBId; // @[Core_1.scala 559:30]
  assign lsuStage_1_io_cache_read_req_ready = dcache_io_read_req_ready; // @[Core_1.scala 572:30]
  assign lsuStage_1_io_cache_read_resp_valid = dcache_io_read_resp_valid; // @[Core_1.scala 572:30]
  assign lsuStage_1_io_cache_read_resp_bits_data = dcache_io_read_resp_bits_data; // @[Core_1.scala 572:30]
  assign lsuStage_1_io_cache_write_req_ready = dcache_io_write_req_ready; // @[Core_1.scala 573:31]
  assign lsuStage_1_io_cache_write_resp_valid = dcache_io_write_resp_valid; // @[Core_1.scala 573:31]
  assign lsuStage_1_io_rob_bits_id = rob_io_deq_bits_id; // @[Core_1.scala 567:31]
  assign lsuStage_1_io_flush = globalBrTaken | reset; // @[Core_1.scala 562:42]
  assign lsuRS_clock = clock;
  assign lsuRS_reset = reset;
  assign lsuRS_io_enq_valid = issue_instFire & issue_lsuValid; // @[Core_1.scala 549:43]
  assign lsuRS_io_enq_bits_op = {{3'd0}, _rob_io_enq_bits_fuOp_T_3}; // @[Core_1.scala 482:23 489:16]
  assign lsuRS_io_enq_bits_opr1 = _issue_chosenDecodesigs_T_45 | _issue_chosenDecodesigs_T_43; // @[Mux.scala 27:73]
  assign lsuRS_io_enq_bits_opr2 = _issue_chosenDecodesigs_T_38 | _issue_chosenDecodesigs_T_36; // @[Mux.scala 27:73]
  assign lsuRS_io_enq_bits_rs1 = issue_chosenDecodesigs_opr1 == 4'h1 ? rs1 : 5'h0; // @[Core_1.scala 266:24]
  assign lsuRS_io_enq_bits_rs2 = issue_chosenDecodesigs_opr2 == 4'h2 ? rs2 : 5'h0; // @[Core_1.scala 267:24]
  assign lsuRS_io_enq_bits_ROBId = {{5'd0}, rob_io_id}; // @[Core_1.scala 482:23 483:19]
  assign lsuRS_io_enq_bits_rs1ROBId = 5'h1f == issue_rs1 ? rob_io_regStatus_31_owner : _GEN_106; // @[Core_1.scala 500:{22,22}]
  assign lsuRS_io_enq_bits_rs2ROBId = 5'h1f == issue_rs1 ? rob_io_regStatus_31_owner : _GEN_106; // @[Core_1.scala 500:{22,22}]
  assign lsuRS_io_enq_bits_immSrc = _issue_chosenDecodesigs_T_31 | _issue_chosenDecodesigs_T_29; // @[Mux.scala 27:73]
  assign lsuRS_io_enq_bits_immSign = _issue_chosenDecodesigs_T[0] & issue_decodeSigs_0_immSign |
    _issue_chosenDecodesigs_T[1] & issue_decodeSigs_1_immSign | _issue_chosenDecodesigs_T[2] &
    issue_decodeSigs_2_immSign | _issue_chosenDecodesigs_T[3] & issue_decodeSigs_3_immSign; // @[Mux.scala 27:73]
  assign lsuRS_io_enq_bits_excpType = _issue_chosenDecodesigs_T_10 | _issue_chosenDecodesigs_T_8; // @[Mux.scala 27:73]
  assign lsuRS_io_enq_bits_pc = issue_stagePc; // @[Core_1.scala 482:23 488:16]
  assign lsuRS_io_enq_bits_inst = _issue_chosenInst_T_10 | _issue_chosenInst_T_8; // @[Mux.scala 27:73]
  assign lsuRS_io_deq_ready = lsuStage_1_io_in_ready; // @[Core_1.scala 553:24]
  assign lsuRS_io_robRead_0_busy = rob_io_read_0_busy; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_0_state = rob_io_read_0_state; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_0_rd = rob_io_read_0_rd; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_0_data = rob_io_read_0_data; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_1_busy = rob_io_read_1_busy; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_1_state = rob_io_read_1_state; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_1_rd = rob_io_read_1_rd; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_1_data = rob_io_read_1_data; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_2_busy = rob_io_read_2_busy; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_2_state = rob_io_read_2_state; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_2_rd = rob_io_read_2_rd; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_2_data = rob_io_read_2_data; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_3_busy = rob_io_read_3_busy; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_3_state = rob_io_read_3_state; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_3_rd = rob_io_read_3_rd; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_3_data = rob_io_read_3_data; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_4_busy = rob_io_read_4_busy; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_4_state = rob_io_read_4_state; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_4_rd = rob_io_read_4_rd; // @[Core_1.scala 646:16]
  assign lsuRS_io_robRead_4_data = rob_io_read_4_data; // @[Core_1.scala 646:16]
  assign lsuRS_io_regStatus_0_owner = rob_io_regStatus_0_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_1_owner = rob_io_regStatus_1_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_2_owner = rob_io_regStatus_2_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_3_owner = rob_io_regStatus_3_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_4_owner = rob_io_regStatus_4_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_5_owner = rob_io_regStatus_5_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_6_owner = rob_io_regStatus_6_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_7_owner = rob_io_regStatus_7_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_8_owner = rob_io_regStatus_8_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_9_owner = rob_io_regStatus_9_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_10_owner = rob_io_regStatus_10_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_11_owner = rob_io_regStatus_11_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_12_owner = rob_io_regStatus_12_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_13_owner = rob_io_regStatus_13_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_14_owner = rob_io_regStatus_14_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_15_owner = rob_io_regStatus_15_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_16_owner = rob_io_regStatus_16_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_17_owner = rob_io_regStatus_17_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_18_owner = rob_io_regStatus_18_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_19_owner = rob_io_regStatus_19_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_20_owner = rob_io_regStatus_20_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_21_owner = rob_io_regStatus_21_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_22_owner = rob_io_regStatus_22_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_23_owner = rob_io_regStatus_23_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_24_owner = rob_io_regStatus_24_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_25_owner = rob_io_regStatus_25_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_26_owner = rob_io_regStatus_26_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_27_owner = rob_io_regStatus_27_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_28_owner = rob_io_regStatus_28_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_29_owner = rob_io_regStatus_29_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_30_owner = rob_io_regStatus_30_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_regStatus_31_owner = rob_io_regStatus_31_owner; // @[Core_1.scala 551:24]
  assign lsuRS_io_cdb_0_valid = aluStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign lsuRS_io_cdb_0_bits_data = aluStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign lsuRS_io_cdb_0_bits_id = aluStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign lsuRS_io_cdb_0_bits_rd = aluStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign lsuRS_io_cdb_1_valid = bruStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign lsuRS_io_cdb_1_bits_data = bruStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign lsuRS_io_cdb_1_bits_id = bruStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign lsuRS_io_cdb_1_bits_rd = bruStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign lsuRS_io_cdb_2_valid = lsuStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign lsuRS_io_cdb_2_bits_data = lsuStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign lsuRS_io_cdb_2_bits_id = lsuStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign lsuRS_io_cdb_2_bits_rd = lsuStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign lsuRS_io_cdb_3_valid = csrStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign lsuRS_io_cdb_3_bits_data = csrStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign lsuRS_io_cdb_3_bits_id = csrStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign lsuRS_io_cdb_3_bits_rd = csrStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign lsuRS_io_rf_0_data = rf_io_r_4_data; // @[Core_1.scala 655:20]
  assign lsuRS_io_rf_1_data = rf_io_r_5_data; // @[Core_1.scala 656:20]
  assign lsuRS_io_flush = globalBrTaken | reset; // @[Core_1.scala 552:37]
  assign csrStage_1_clock = clock;
  assign csrStage_1_reset = reset;
  assign csrStage_1_io_in_valid = csrRS_io_deq_valid; // @[Core_1.scala 583:28]
  assign csrStage_1_io_in_bits_csrOp = csrRS_io_deq_bits_op[2:0]; // @[Core_1.scala 585:33]
  assign csrStage_1_io_in_bits_excpType = csrRS_io_deq_bits_excpType; // @[Core_1.scala 584:36]
  assign csrStage_1_io_in_bits_rs1Val = csrRS_io_deq_bits_rs1Val; // @[Core_1.scala 588:34]
  assign csrStage_1_io_in_bits_inst = csrRS_io_deq_bits_inst; // @[Core_1.scala 586:32]
  assign csrStage_1_io_in_bits_id = csrRS_io_deq_bits_ROBId; // @[Core_1.scala 587:30]
  assign csrStage_1_io_flush = globalBrTaken | reset; // @[Core_1.scala 590:42]
  assign csrRS_clock = clock;
  assign csrRS_reset = reset;
  assign csrRS_io_enq_valid = issue_instFire & issue_csrValid; // @[Core_1.scala 577:43]
  assign csrRS_io_enq_bits_op = {{3'd0}, _rob_io_enq_bits_fuOp_T_3}; // @[Core_1.scala 482:23 489:16]
  assign csrRS_io_enq_bits_opr1 = _issue_chosenDecodesigs_T_45 | _issue_chosenDecodesigs_T_43; // @[Mux.scala 27:73]
  assign csrRS_io_enq_bits_opr2 = _issue_chosenDecodesigs_T_38 | _issue_chosenDecodesigs_T_36; // @[Mux.scala 27:73]
  assign csrRS_io_enq_bits_rs1 = issue_chosenDecodesigs_opr1 == 4'h1 ? rs1 : 5'h0; // @[Core_1.scala 266:24]
  assign csrRS_io_enq_bits_rs2 = issue_chosenDecodesigs_opr2 == 4'h2 ? rs2 : 5'h0; // @[Core_1.scala 267:24]
  assign csrRS_io_enq_bits_ROBId = {{5'd0}, rob_io_id}; // @[Core_1.scala 482:23 483:19]
  assign csrRS_io_enq_bits_rs1ROBId = 5'h1f == issue_rs1 ? rob_io_regStatus_31_owner : _GEN_106; // @[Core_1.scala 500:{22,22}]
  assign csrRS_io_enq_bits_rs2ROBId = 5'h1f == issue_rs1 ? rob_io_regStatus_31_owner : _GEN_106; // @[Core_1.scala 500:{22,22}]
  assign csrRS_io_enq_bits_immSrc = _issue_chosenDecodesigs_T_31 | _issue_chosenDecodesigs_T_29; // @[Mux.scala 27:73]
  assign csrRS_io_enq_bits_immSign = _issue_chosenDecodesigs_T[0] & issue_decodeSigs_0_immSign |
    _issue_chosenDecodesigs_T[1] & issue_decodeSigs_1_immSign | _issue_chosenDecodesigs_T[2] &
    issue_decodeSigs_2_immSign | _issue_chosenDecodesigs_T[3] & issue_decodeSigs_3_immSign; // @[Mux.scala 27:73]
  assign csrRS_io_enq_bits_excpType = _issue_chosenDecodesigs_T_10 | _issue_chosenDecodesigs_T_8; // @[Mux.scala 27:73]
  assign csrRS_io_enq_bits_pc = issue_stagePc; // @[Core_1.scala 482:23 488:16]
  assign csrRS_io_enq_bits_inst = _issue_chosenInst_T_10 | _issue_chosenInst_T_8; // @[Mux.scala 27:73]
  assign csrRS_io_deq_ready = csrStage_1_io_in_ready; // @[Core_1.scala 581:24]
  assign csrRS_io_robRead_0_busy = rob_io_read_0_busy; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_0_state = rob_io_read_0_state; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_0_rd = rob_io_read_0_rd; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_0_data = rob_io_read_0_data; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_1_busy = rob_io_read_1_busy; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_1_state = rob_io_read_1_state; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_1_rd = rob_io_read_1_rd; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_1_data = rob_io_read_1_data; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_2_busy = rob_io_read_2_busy; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_2_state = rob_io_read_2_state; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_2_rd = rob_io_read_2_rd; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_2_data = rob_io_read_2_data; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_3_busy = rob_io_read_3_busy; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_3_state = rob_io_read_3_state; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_3_rd = rob_io_read_3_rd; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_3_data = rob_io_read_3_data; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_4_busy = rob_io_read_4_busy; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_4_state = rob_io_read_4_state; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_4_rd = rob_io_read_4_rd; // @[Core_1.scala 646:16]
  assign csrRS_io_robRead_4_data = rob_io_read_4_data; // @[Core_1.scala 646:16]
  assign csrRS_io_regStatus_0_owner = rob_io_regStatus_0_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_1_owner = rob_io_regStatus_1_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_2_owner = rob_io_regStatus_2_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_3_owner = rob_io_regStatus_3_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_4_owner = rob_io_regStatus_4_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_5_owner = rob_io_regStatus_5_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_6_owner = rob_io_regStatus_6_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_7_owner = rob_io_regStatus_7_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_8_owner = rob_io_regStatus_8_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_9_owner = rob_io_regStatus_9_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_10_owner = rob_io_regStatus_10_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_11_owner = rob_io_regStatus_11_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_12_owner = rob_io_regStatus_12_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_13_owner = rob_io_regStatus_13_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_14_owner = rob_io_regStatus_14_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_15_owner = rob_io_regStatus_15_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_16_owner = rob_io_regStatus_16_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_17_owner = rob_io_regStatus_17_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_18_owner = rob_io_regStatus_18_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_19_owner = rob_io_regStatus_19_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_20_owner = rob_io_regStatus_20_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_21_owner = rob_io_regStatus_21_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_22_owner = rob_io_regStatus_22_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_23_owner = rob_io_regStatus_23_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_24_owner = rob_io_regStatus_24_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_25_owner = rob_io_regStatus_25_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_26_owner = rob_io_regStatus_26_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_27_owner = rob_io_regStatus_27_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_28_owner = rob_io_regStatus_28_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_29_owner = rob_io_regStatus_29_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_30_owner = rob_io_regStatus_30_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_regStatus_31_owner = rob_io_regStatus_31_owner; // @[Core_1.scala 579:24]
  assign csrRS_io_cdb_0_valid = aluStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign csrRS_io_cdb_0_bits_data = aluStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign csrRS_io_cdb_0_bits_id = aluStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign csrRS_io_cdb_0_bits_rd = aluStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign csrRS_io_cdb_1_valid = bruStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign csrRS_io_cdb_1_bits_data = bruStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign csrRS_io_cdb_1_bits_id = bruStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign csrRS_io_cdb_1_bits_rd = bruStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign csrRS_io_cdb_2_valid = lsuStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign csrRS_io_cdb_2_bits_data = lsuStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign csrRS_io_cdb_2_bits_id = lsuStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign csrRS_io_cdb_2_bits_rd = lsuStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign csrRS_io_cdb_3_valid = csrStage_1_io_out_valid; // @[Core_1.scala 634:21]
  assign csrRS_io_cdb_3_bits_data = csrStage_1_io_out_bits_data; // @[Core_1.scala 635:25]
  assign csrRS_io_cdb_3_bits_id = csrStage_1_io_out_bits_id; // @[Core_1.scala 637:23]
  assign csrRS_io_cdb_3_bits_rd = csrStage_1_io_out_bits_rd; // @[Core_1.scala 636:23]
  assign csrRS_io_rf_0_data = rf_io_r_6_data; // @[Core_1.scala 657:20]
  assign csrRS_io_rf_1_data = rf_io_r_7_data; // @[Core_1.scala 658:20]
  assign csrRS_io_flush = globalBrTaken | reset; // @[Core_1.scala 580:37]
  assign edgeBackPressure_clock = clock;
  assign edgeBackPressure_io_in = ib_io_status_back_pressure; // @[Core_1.scala 131:28]
  assign fetch_pendingBranch_clock = clock;
  assign fetch_pendingBranch_reset = reset;
  assign fetch_pendingBranch_io_enq_valid = globalBrTaken; // @[Core_1.scala 137:38]
  assign fetch_pendingBranch_io_enq_bits = csrExcpValid ? csrExcpAddr : bruBrAddr; // @[Core_1.scala 105:27]
  assign fetch_pendingBranch_io_deq_ready = icache_io_read_req_ready; // @[Core_1.scala 138:38]
  assign dec_decoders_0_io_inst = dec_inst_0_inst; // @[Core_1.scala 201:33]
  assign dec_decoders_1_io_inst = dec_inst_1_inst; // @[Core_1.scala 201:33]
  assign dec_decoders_2_io_inst = dec_inst_2_inst; // @[Core_1.scala 201:33]
  assign dec_decoders_3_io_inst = dec_inst_3_inst; // @[Core_1.scala 201:33]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_read_req_valid = lsuStage_1_io_cache_read_req_valid; // @[Core_1.scala 572:30]
  assign dcache_io_read_req_bits_addr = lsuStage_1_io_cache_read_req_bits_addr; // @[Core_1.scala 572:30]
  assign dcache_io_read_resp_ready = lsuStage_1_io_cache_read_resp_ready; // @[Core_1.scala 572:30]
  assign dcache_io_write_req_valid = lsuStage_1_io_cache_write_req_valid; // @[Core_1.scala 573:31]
  assign dcache_io_write_req_bits_addr = lsuStage_1_io_cache_write_req_bits_addr; // @[Core_1.scala 573:31]
  assign dcache_io_write_req_bits_data = lsuStage_1_io_cache_write_req_bits_data; // @[Core_1.scala 573:31]
  assign dcache_io_write_req_bits_mask = lsuStage_1_io_cache_write_req_bits_mask; // @[Core_1.scala 573:31]
  assign dcache_io_write_resp_ready = lsuStage_1_io_cache_write_resp_ready; // @[Core_1.scala 573:31]
  assign dcache_io_tlbus_req_ready = xbar_io_masterFace_in_1_ready; // @[Core_1.scala 701:25]
  assign dcache_io_tlbus_resp_valid = xbar_io_masterFace_out_1_valid; // @[Core_1.scala 702:26]
  assign dcache_io_tlbus_resp_bits_opcode = xbar_io_masterFace_out_1_bits_opcode; // @[Core_1.scala 702:26]
  assign dcache_io_tlbus_resp_bits_data = xbar_io_masterFace_out_1_bits_data; // @[Core_1.scala 702:26]
  assign dcache_io_flush = globalBrTaken; // @[Core_1.scala 571:21]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_masterFace_in_0_valid = icache_io_tlbus_req_valid; // @[Core_1.scala 698:25]
  assign xbar_io_masterFace_in_0_bits_address = icache_io_tlbus_req_bits_address; // @[Core_1.scala 698:25]
  assign xbar_io_masterFace_in_1_valid = dcache_io_tlbus_req_valid; // @[Core_1.scala 701:25]
  assign xbar_io_masterFace_in_1_bits_opcode = dcache_io_tlbus_req_bits_opcode; // @[Core_1.scala 701:25]
  assign xbar_io_masterFace_in_1_bits_address = dcache_io_tlbus_req_bits_address; // @[Core_1.scala 701:25]
  assign xbar_io_masterFace_in_1_bits_data = dcache_io_tlbus_req_bits_data; // @[Core_1.scala 701:25]
  assign xbar_io_slaveFace_in_0_ready = rom_io_req_ready; // @[Core_1.scala 704:16]
  assign xbar_io_slaveFace_out_0_valid = rom_io_resp_valid; // @[Core_1.scala 705:17]
  assign xbar_io_slaveFace_out_0_bits_opcode = rom_io_resp_bits_opcode; // @[Core_1.scala 705:17]
  assign xbar_io_slaveFace_out_0_bits_data = rom_io_resp_bits_data; // @[Core_1.scala 705:17]
  assign rom_clock = clock;
  assign rom_reset = reset;
  assign rom_io_req_valid = xbar_io_slaveFace_in_0_valid; // @[Core_1.scala 704:16]
  assign rom_io_req_bits_opcode = xbar_io_slaveFace_in_0_bits_opcode; // @[Core_1.scala 704:16]
  assign rom_io_req_bits_size = xbar_io_slaveFace_in_0_bits_size; // @[Core_1.scala 704:16]
  assign rom_io_req_bits_address = xbar_io_slaveFace_in_0_bits_address; // @[Core_1.scala 704:16]
  assign rom_io_req_bits_data = xbar_io_slaveFace_in_0_bits_data; // @[Core_1.scala 704:16]
  assign rom_io_resp_ready = xbar_io_slaveFace_out_0_ready; // @[Core_1.scala 705:17]
  always @(posedge clock) begin
    if (reset) begin // @[Core_1.scala 114:24]
      pcReg <= 32'h0; // @[Core_1.scala 114:24]
    end else if (_lastPc_T & _preFetchInst_T_2) begin // @[Core_1.scala 156:49]
      if (brTaken) begin // @[Core_1.scala 159:18]
        pcReg <= fetch_pendingBranch_io_deq_bits;
      end else if (isAlignAddr) begin // @[Core_1.scala 119:22]
        pcReg <= _pcNext4_T_1;
      end else begin
        pcReg <= _pcNext4_T_8;
      end
    end
    if (_lastPc_T) begin // @[Reg.scala 20:18]
      lastPc <= icache_io_read_req_bits_addr; // @[Reg.scala 20:22]
    end
    firstFire <= reset | _GEN_3; // @[Reg.scala 35:{20,20}]
    if (globalBrTaken) begin // @[Reg.scala 20:18]
      if (csrExcpValid) begin // @[Core_1.scala 105:27]
        blockAddr <= csrExcpAddr;
      end else begin
        blockAddr <= bruBrAddr;
      end
    end
    if (reset) begin // @[Core_1.scala 166:29]
      blockValid <= 1'h0; // @[Core_1.scala 166:29]
    end else begin
      blockValid <= _GEN_7;
    end
    if (reset) begin // @[Core_1.scala 186:27]
      dec_full <= 1'h0; // @[Core_1.scala 186:27]
    end else if (_ib_io_in_bits_flush_T_1) begin // @[Core_1.scala 212:21]
      dec_full <= 1'h0; // @[Core_1.scala 213:18]
    end else begin
      dec_full <= _GEN_18;
    end
    if (reset) begin // @[Core_1.scala 224:29]
      issue_full <= 1'h0; // @[Core_1.scala 224:29]
    end else if (_ib_io_in_bits_flush_T_1) begin // @[Core_1.scala 257:23]
      issue_full <= 1'h0; // @[Core_1.scala 258:20]
    end else begin
      issue_full <= _GEN_71;
    end
    if (reset) begin // @[Core_1.scala 231:28]
      issue_ptr <= 2'h0; // @[Core_1.scala 231:28]
    end else if (_ib_io_in_bits_flush_T_1) begin // @[Core_1.scala 257:23]
      issue_ptr <= 2'h0; // @[Core_1.scala 259:19]
    end else if (issue_fire) begin // @[Core_1.scala 248:22]
      issue_ptr <= 2'h0; // @[Core_1.scala 248:34]
    end else if (issue_instFire) begin // @[Core_1.scala 249:31]
      issue_ptr <= _issue_ptr_T_1; // @[Core_1.scala 249:43]
    end
    if (dec_fire) begin // @[Reg.scala 20:18]
      issue_instValid <= _issue_instValid_T; // @[Reg.scala 20:22]
    end
    if (dec_latch) begin // @[Reg.scala 20:18]
      dec_inst_0_inst <= ib_io_out_bits_inst_0_inst; // @[Reg.scala 20:22]
    end
    if (_ib_io_in_bits_flush_T_1) begin // @[Core_1.scala 212:21]
      dec_inst_0_valid <= 1'h0; // @[Core_1.scala 214:40]
    end else if (dec_latch) begin // @[Reg.scala 20:18]
      dec_inst_0_valid <= ib_io_out_bits_inst_0_valid; // @[Reg.scala 20:22]
    end
    if (dec_latch) begin // @[Reg.scala 20:18]
      dec_inst_1_inst <= ib_io_out_bits_inst_1_inst; // @[Reg.scala 20:22]
    end
    if (_ib_io_in_bits_flush_T_1) begin // @[Core_1.scala 212:21]
      dec_inst_1_valid <= 1'h0; // @[Core_1.scala 214:40]
    end else if (dec_latch) begin // @[Reg.scala 20:18]
      dec_inst_1_valid <= ib_io_out_bits_inst_1_valid; // @[Reg.scala 20:22]
    end
    if (dec_latch) begin // @[Reg.scala 20:18]
      dec_inst_2_inst <= ib_io_out_bits_inst_2_inst; // @[Reg.scala 20:22]
    end
    if (_ib_io_in_bits_flush_T_1) begin // @[Core_1.scala 212:21]
      dec_inst_2_valid <= 1'h0; // @[Core_1.scala 214:40]
    end else if (dec_latch) begin // @[Reg.scala 20:18]
      dec_inst_2_valid <= ib_io_out_bits_inst_2_valid; // @[Reg.scala 20:22]
    end
    if (dec_latch) begin // @[Reg.scala 20:18]
      dec_inst_3_inst <= ib_io_out_bits_inst_3_inst; // @[Reg.scala 20:22]
    end
    if (_ib_io_in_bits_flush_T_1) begin // @[Core_1.scala 212:21]
      dec_inst_3_valid <= 1'h0; // @[Core_1.scala 214:40]
    end else if (dec_latch) begin // @[Reg.scala 20:18]
      dec_inst_3_valid <= ib_io_out_bits_inst_3_valid; // @[Reg.scala 20:22]
    end
    if (dec_latch) begin // @[Reg.scala 20:18]
      dec_pc <= ib_io_out_bits_pc; // @[Reg.scala 20:22]
    end
    if (dec_fire) begin // @[Reg.scala 20:18]
      issue_pc <= dec_pc; // @[Reg.scala 20:22]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_0_brType <= dec_decodeSigs_0_brType; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_0_lsuOp <= dec_decodeSigs_0_lsuOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_0_aluOp <= dec_decodeSigs_0_aluOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_0_opr1 <= dec_decodeSigs_0_opr1; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_0_opr2 <= dec_decodeSigs_0_opr2; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_0_immSrc <= dec_decodeSigs_0_immSrc; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_0_immSign <= dec_decodeSigs_0_immSign; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_0_csrOp <= dec_decodeSigs_0_csrOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_0_excpType <= dec_decodeSigs_0_excpType; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_1_brType <= dec_decodeSigs_1_brType; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_1_lsuOp <= dec_decodeSigs_1_lsuOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_1_aluOp <= dec_decodeSigs_1_aluOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_1_opr1 <= dec_decodeSigs_1_opr1; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_1_opr2 <= dec_decodeSigs_1_opr2; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_1_immSrc <= dec_decodeSigs_1_immSrc; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_1_immSign <= dec_decodeSigs_1_immSign; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_1_csrOp <= dec_decodeSigs_1_csrOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_1_excpType <= dec_decodeSigs_1_excpType; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_2_brType <= dec_decodeSigs_2_brType; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_2_lsuOp <= dec_decodeSigs_2_lsuOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_2_aluOp <= dec_decodeSigs_2_aluOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_2_opr1 <= dec_decodeSigs_2_opr1; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_2_opr2 <= dec_decodeSigs_2_opr2; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_2_immSrc <= dec_decodeSigs_2_immSrc; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_2_immSign <= dec_decodeSigs_2_immSign; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_2_csrOp <= dec_decodeSigs_2_csrOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_2_excpType <= dec_decodeSigs_2_excpType; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_3_brType <= dec_decodeSigs_3_brType; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_3_lsuOp <= dec_decodeSigs_3_lsuOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_3_aluOp <= dec_decodeSigs_3_aluOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_3_opr1 <= dec_decodeSigs_3_opr1; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_3_opr2 <= dec_decodeSigs_3_opr2; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_3_immSrc <= dec_decodeSigs_3_immSrc; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_3_immSign <= dec_decodeSigs_3_immSign; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_3_csrOp <= dec_decodeSigs_3_csrOp; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_decodeSigs_3_excpType <= dec_decodeSigs_3_excpType; // @[Core_1.scala 235:33]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_inst_0 <= dec_inst_0_inst; // @[Core_1.scala 236:27]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_inst_1 <= dec_inst_1_inst; // @[Core_1.scala 236:27]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_inst_2 <= dec_inst_2_inst; // @[Core_1.scala 236:27]
    end
    if (dec_fire) begin // @[Core_1.scala 234:27]
      issue_inst_3 <= dec_inst_3_inst; // @[Core_1.scala 236:27]
    end
    io_out_state_instState_REG_commit <= rob_io_deq_ready & rob_io_deq_valid; // @[Decoupled.scala 51:35]
    io_out_state_instState_REG_pc <= rob_io_deq_bits_pc; // @[Core_1.scala 673:25 676:18]
    io_out_state_instState_REG_inst <= rob_io_deq_bits_inst; // @[Core_1.scala 673:25 675:20]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_12 <= 3'h1 & issue_full | _issue_ready_T)) begin
          $fwrite(32'h80000002,
            "Assertion failed: more than one op valid! %d %d %d %d inst=> %x aluOp=> %d bruOp=> %d lsuOp=> %d csrOp=> %d excpType=> %d\n    at Core_1.scala:276 assert(((PopCount(VecInit(Seq(issue_aluValid, issue_bruValid, issue_lsuValid, issue_csrValid))) <= 1.U && issue_full) || !issue_full),\n"
            ,issue_aluValid,issue_bruValid,issue_lsuValid,issue_csrValid,issue_chosenInst,issue_chosenDecodesigs_aluOp,
            issue_chosenDecodesigs_brType,issue_chosenDecodesigs_lsuOp,issue_chosenDecodesigs_csrOp,
            issue_chosenDecodesigs_excpType); // @[Core_1.scala 276:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_12 <= 3'h1 & issue_full | _issue_ready_T) & ~reset) begin
          $fatal; // @[Core_1.scala 276:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  lastPc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  firstFire = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  blockAddr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  blockValid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dec_full = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  issue_full = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  issue_ptr = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  issue_instValid = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  dec_inst_0_inst = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  dec_inst_0_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dec_inst_1_inst = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  dec_inst_1_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  dec_inst_2_inst = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  dec_inst_2_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  dec_inst_3_inst = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  dec_inst_3_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  dec_pc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  issue_pc = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  issue_decodeSigs_0_brType = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  issue_decodeSigs_0_lsuOp = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  issue_decodeSigs_0_aluOp = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  issue_decodeSigs_0_opr1 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  issue_decodeSigs_0_opr2 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  issue_decodeSigs_0_immSrc = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  issue_decodeSigs_0_immSign = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  issue_decodeSigs_0_csrOp = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  issue_decodeSigs_0_excpType = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  issue_decodeSigs_1_brType = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  issue_decodeSigs_1_lsuOp = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  issue_decodeSigs_1_aluOp = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  issue_decodeSigs_1_opr1 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  issue_decodeSigs_1_opr2 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  issue_decodeSigs_1_immSrc = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  issue_decodeSigs_1_immSign = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  issue_decodeSigs_1_csrOp = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  issue_decodeSigs_1_excpType = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  issue_decodeSigs_2_brType = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  issue_decodeSigs_2_lsuOp = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  issue_decodeSigs_2_aluOp = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  issue_decodeSigs_2_opr1 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  issue_decodeSigs_2_opr2 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  issue_decodeSigs_2_immSrc = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  issue_decodeSigs_2_immSign = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  issue_decodeSigs_2_csrOp = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  issue_decodeSigs_2_excpType = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  issue_decodeSigs_3_brType = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  issue_decodeSigs_3_lsuOp = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  issue_decodeSigs_3_aluOp = _RAND_48[4:0];
  _RAND_49 = {1{`RANDOM}};
  issue_decodeSigs_3_opr1 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  issue_decodeSigs_3_opr2 = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  issue_decodeSigs_3_immSrc = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  issue_decodeSigs_3_immSign = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  issue_decodeSigs_3_csrOp = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  issue_decodeSigs_3_excpType = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  issue_inst_0 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  issue_inst_1 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  issue_inst_2 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  issue_inst_3 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  io_out_state_instState_REG_commit = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  io_out_state_instState_REG_pc = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  io_out_state_instState_REG_inst = _RAND_61[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
