module BankRAM_2P_112(
  input         clock,
  input         reset,
  input  [7:0]  io_r_addr,
  output [19:0] io_r_data,
  input         io_w_en,
  input  [7:0]  io_w_addr,
  input  [19:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] mem [0:255]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_129_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_130_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_131_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_132_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_133_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_134_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_135_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_136_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_137_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_138_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_139_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_140_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_141_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_142_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_143_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_144_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_145_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_146_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_147_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_148_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_149_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_150_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_151_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_152_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_153_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_154_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_155_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_156_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_157_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_158_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_159_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_160_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_161_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_162_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_163_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_164_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_165_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_166_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_167_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_168_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_169_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_170_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_171_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_172_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_173_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_174_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_175_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_176_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_177_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_178_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_179_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_180_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_181_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_182_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_183_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_184_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_185_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_186_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_187_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_188_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_189_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_190_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_191_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_192_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_193_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_194_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_195_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_196_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_197_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_198_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_199_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_200_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_201_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_202_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_203_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_204_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_205_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_206_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_207_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_208_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_209_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_210_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_211_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_212_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_213_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_214_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_215_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_216_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_217_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_218_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_219_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_220_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_221_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_222_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_223_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_224_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_225_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_226_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_227_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_228_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_229_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_230_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_231_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_232_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_233_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_234_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_235_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_236_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_237_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_238_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_239_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_240_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_241_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_242_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_243_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_244_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_245_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_246_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_247_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_248_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_249_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_250_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_251_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_252_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_253_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_254_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_255_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_256_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [7:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 20'h0;
  assign mem_MPORT_addr = 8'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 20'h0;
  assign mem_MPORT_1_addr = 8'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 20'h0;
  assign mem_MPORT_2_addr = 8'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 20'h0;
  assign mem_MPORT_3_addr = 8'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 20'h0;
  assign mem_MPORT_4_addr = 8'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 20'h0;
  assign mem_MPORT_5_addr = 8'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 20'h0;
  assign mem_MPORT_6_addr = 8'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 20'h0;
  assign mem_MPORT_7_addr = 8'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 20'h0;
  assign mem_MPORT_8_addr = 8'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 20'h0;
  assign mem_MPORT_9_addr = 8'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 20'h0;
  assign mem_MPORT_10_addr = 8'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 20'h0;
  assign mem_MPORT_11_addr = 8'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 20'h0;
  assign mem_MPORT_12_addr = 8'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 20'h0;
  assign mem_MPORT_13_addr = 8'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 20'h0;
  assign mem_MPORT_14_addr = 8'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 20'h0;
  assign mem_MPORT_15_addr = 8'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 20'h0;
  assign mem_MPORT_16_addr = 8'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 20'h0;
  assign mem_MPORT_17_addr = 8'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 20'h0;
  assign mem_MPORT_18_addr = 8'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 20'h0;
  assign mem_MPORT_19_addr = 8'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 20'h0;
  assign mem_MPORT_20_addr = 8'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 20'h0;
  assign mem_MPORT_21_addr = 8'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 20'h0;
  assign mem_MPORT_22_addr = 8'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 20'h0;
  assign mem_MPORT_23_addr = 8'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 20'h0;
  assign mem_MPORT_24_addr = 8'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 20'h0;
  assign mem_MPORT_25_addr = 8'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 20'h0;
  assign mem_MPORT_26_addr = 8'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 20'h0;
  assign mem_MPORT_27_addr = 8'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 20'h0;
  assign mem_MPORT_28_addr = 8'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 20'h0;
  assign mem_MPORT_29_addr = 8'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 20'h0;
  assign mem_MPORT_30_addr = 8'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 20'h0;
  assign mem_MPORT_31_addr = 8'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 20'h0;
  assign mem_MPORT_32_addr = 8'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 20'h0;
  assign mem_MPORT_33_addr = 8'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 20'h0;
  assign mem_MPORT_34_addr = 8'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 20'h0;
  assign mem_MPORT_35_addr = 8'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 20'h0;
  assign mem_MPORT_36_addr = 8'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 20'h0;
  assign mem_MPORT_37_addr = 8'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 20'h0;
  assign mem_MPORT_38_addr = 8'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 20'h0;
  assign mem_MPORT_39_addr = 8'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 20'h0;
  assign mem_MPORT_40_addr = 8'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 20'h0;
  assign mem_MPORT_41_addr = 8'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 20'h0;
  assign mem_MPORT_42_addr = 8'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 20'h0;
  assign mem_MPORT_43_addr = 8'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 20'h0;
  assign mem_MPORT_44_addr = 8'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 20'h0;
  assign mem_MPORT_45_addr = 8'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 20'h0;
  assign mem_MPORT_46_addr = 8'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 20'h0;
  assign mem_MPORT_47_addr = 8'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 20'h0;
  assign mem_MPORT_48_addr = 8'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 20'h0;
  assign mem_MPORT_49_addr = 8'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 20'h0;
  assign mem_MPORT_50_addr = 8'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 20'h0;
  assign mem_MPORT_51_addr = 8'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 20'h0;
  assign mem_MPORT_52_addr = 8'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 20'h0;
  assign mem_MPORT_53_addr = 8'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 20'h0;
  assign mem_MPORT_54_addr = 8'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 20'h0;
  assign mem_MPORT_55_addr = 8'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 20'h0;
  assign mem_MPORT_56_addr = 8'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 20'h0;
  assign mem_MPORT_57_addr = 8'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 20'h0;
  assign mem_MPORT_58_addr = 8'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 20'h0;
  assign mem_MPORT_59_addr = 8'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 20'h0;
  assign mem_MPORT_60_addr = 8'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 20'h0;
  assign mem_MPORT_61_addr = 8'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 20'h0;
  assign mem_MPORT_62_addr = 8'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 20'h0;
  assign mem_MPORT_63_addr = 8'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 20'h0;
  assign mem_MPORT_64_addr = 8'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 20'h0;
  assign mem_MPORT_65_addr = 8'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 20'h0;
  assign mem_MPORT_66_addr = 8'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 20'h0;
  assign mem_MPORT_67_addr = 8'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 20'h0;
  assign mem_MPORT_68_addr = 8'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 20'h0;
  assign mem_MPORT_69_addr = 8'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 20'h0;
  assign mem_MPORT_70_addr = 8'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 20'h0;
  assign mem_MPORT_71_addr = 8'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 20'h0;
  assign mem_MPORT_72_addr = 8'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 20'h0;
  assign mem_MPORT_73_addr = 8'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 20'h0;
  assign mem_MPORT_74_addr = 8'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 20'h0;
  assign mem_MPORT_75_addr = 8'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 20'h0;
  assign mem_MPORT_76_addr = 8'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 20'h0;
  assign mem_MPORT_77_addr = 8'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 20'h0;
  assign mem_MPORT_78_addr = 8'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 20'h0;
  assign mem_MPORT_79_addr = 8'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 20'h0;
  assign mem_MPORT_80_addr = 8'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 20'h0;
  assign mem_MPORT_81_addr = 8'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 20'h0;
  assign mem_MPORT_82_addr = 8'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 20'h0;
  assign mem_MPORT_83_addr = 8'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 20'h0;
  assign mem_MPORT_84_addr = 8'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 20'h0;
  assign mem_MPORT_85_addr = 8'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 20'h0;
  assign mem_MPORT_86_addr = 8'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 20'h0;
  assign mem_MPORT_87_addr = 8'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 20'h0;
  assign mem_MPORT_88_addr = 8'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 20'h0;
  assign mem_MPORT_89_addr = 8'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 20'h0;
  assign mem_MPORT_90_addr = 8'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 20'h0;
  assign mem_MPORT_91_addr = 8'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 20'h0;
  assign mem_MPORT_92_addr = 8'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 20'h0;
  assign mem_MPORT_93_addr = 8'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 20'h0;
  assign mem_MPORT_94_addr = 8'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 20'h0;
  assign mem_MPORT_95_addr = 8'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 20'h0;
  assign mem_MPORT_96_addr = 8'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 20'h0;
  assign mem_MPORT_97_addr = 8'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 20'h0;
  assign mem_MPORT_98_addr = 8'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 20'h0;
  assign mem_MPORT_99_addr = 8'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 20'h0;
  assign mem_MPORT_100_addr = 8'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 20'h0;
  assign mem_MPORT_101_addr = 8'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 20'h0;
  assign mem_MPORT_102_addr = 8'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 20'h0;
  assign mem_MPORT_103_addr = 8'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 20'h0;
  assign mem_MPORT_104_addr = 8'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 20'h0;
  assign mem_MPORT_105_addr = 8'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 20'h0;
  assign mem_MPORT_106_addr = 8'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 20'h0;
  assign mem_MPORT_107_addr = 8'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 20'h0;
  assign mem_MPORT_108_addr = 8'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 20'h0;
  assign mem_MPORT_109_addr = 8'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 20'h0;
  assign mem_MPORT_110_addr = 8'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 20'h0;
  assign mem_MPORT_111_addr = 8'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 20'h0;
  assign mem_MPORT_112_addr = 8'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 20'h0;
  assign mem_MPORT_113_addr = 8'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 20'h0;
  assign mem_MPORT_114_addr = 8'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 20'h0;
  assign mem_MPORT_115_addr = 8'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 20'h0;
  assign mem_MPORT_116_addr = 8'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 20'h0;
  assign mem_MPORT_117_addr = 8'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 20'h0;
  assign mem_MPORT_118_addr = 8'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 20'h0;
  assign mem_MPORT_119_addr = 8'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 20'h0;
  assign mem_MPORT_120_addr = 8'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 20'h0;
  assign mem_MPORT_121_addr = 8'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 20'h0;
  assign mem_MPORT_122_addr = 8'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 20'h0;
  assign mem_MPORT_123_addr = 8'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 20'h0;
  assign mem_MPORT_124_addr = 8'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 20'h0;
  assign mem_MPORT_125_addr = 8'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 20'h0;
  assign mem_MPORT_126_addr = 8'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 20'h0;
  assign mem_MPORT_127_addr = 8'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 20'h0;
  assign mem_MPORT_128_addr = 8'h80;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = reset;
  assign mem_MPORT_129_data = 20'h0;
  assign mem_MPORT_129_addr = 8'h81;
  assign mem_MPORT_129_mask = 1'h1;
  assign mem_MPORT_129_en = reset;
  assign mem_MPORT_130_data = 20'h0;
  assign mem_MPORT_130_addr = 8'h82;
  assign mem_MPORT_130_mask = 1'h1;
  assign mem_MPORT_130_en = reset;
  assign mem_MPORT_131_data = 20'h0;
  assign mem_MPORT_131_addr = 8'h83;
  assign mem_MPORT_131_mask = 1'h1;
  assign mem_MPORT_131_en = reset;
  assign mem_MPORT_132_data = 20'h0;
  assign mem_MPORT_132_addr = 8'h84;
  assign mem_MPORT_132_mask = 1'h1;
  assign mem_MPORT_132_en = reset;
  assign mem_MPORT_133_data = 20'h0;
  assign mem_MPORT_133_addr = 8'h85;
  assign mem_MPORT_133_mask = 1'h1;
  assign mem_MPORT_133_en = reset;
  assign mem_MPORT_134_data = 20'h0;
  assign mem_MPORT_134_addr = 8'h86;
  assign mem_MPORT_134_mask = 1'h1;
  assign mem_MPORT_134_en = reset;
  assign mem_MPORT_135_data = 20'h0;
  assign mem_MPORT_135_addr = 8'h87;
  assign mem_MPORT_135_mask = 1'h1;
  assign mem_MPORT_135_en = reset;
  assign mem_MPORT_136_data = 20'h0;
  assign mem_MPORT_136_addr = 8'h88;
  assign mem_MPORT_136_mask = 1'h1;
  assign mem_MPORT_136_en = reset;
  assign mem_MPORT_137_data = 20'h0;
  assign mem_MPORT_137_addr = 8'h89;
  assign mem_MPORT_137_mask = 1'h1;
  assign mem_MPORT_137_en = reset;
  assign mem_MPORT_138_data = 20'h0;
  assign mem_MPORT_138_addr = 8'h8a;
  assign mem_MPORT_138_mask = 1'h1;
  assign mem_MPORT_138_en = reset;
  assign mem_MPORT_139_data = 20'h0;
  assign mem_MPORT_139_addr = 8'h8b;
  assign mem_MPORT_139_mask = 1'h1;
  assign mem_MPORT_139_en = reset;
  assign mem_MPORT_140_data = 20'h0;
  assign mem_MPORT_140_addr = 8'h8c;
  assign mem_MPORT_140_mask = 1'h1;
  assign mem_MPORT_140_en = reset;
  assign mem_MPORT_141_data = 20'h0;
  assign mem_MPORT_141_addr = 8'h8d;
  assign mem_MPORT_141_mask = 1'h1;
  assign mem_MPORT_141_en = reset;
  assign mem_MPORT_142_data = 20'h0;
  assign mem_MPORT_142_addr = 8'h8e;
  assign mem_MPORT_142_mask = 1'h1;
  assign mem_MPORT_142_en = reset;
  assign mem_MPORT_143_data = 20'h0;
  assign mem_MPORT_143_addr = 8'h8f;
  assign mem_MPORT_143_mask = 1'h1;
  assign mem_MPORT_143_en = reset;
  assign mem_MPORT_144_data = 20'h0;
  assign mem_MPORT_144_addr = 8'h90;
  assign mem_MPORT_144_mask = 1'h1;
  assign mem_MPORT_144_en = reset;
  assign mem_MPORT_145_data = 20'h0;
  assign mem_MPORT_145_addr = 8'h91;
  assign mem_MPORT_145_mask = 1'h1;
  assign mem_MPORT_145_en = reset;
  assign mem_MPORT_146_data = 20'h0;
  assign mem_MPORT_146_addr = 8'h92;
  assign mem_MPORT_146_mask = 1'h1;
  assign mem_MPORT_146_en = reset;
  assign mem_MPORT_147_data = 20'h0;
  assign mem_MPORT_147_addr = 8'h93;
  assign mem_MPORT_147_mask = 1'h1;
  assign mem_MPORT_147_en = reset;
  assign mem_MPORT_148_data = 20'h0;
  assign mem_MPORT_148_addr = 8'h94;
  assign mem_MPORT_148_mask = 1'h1;
  assign mem_MPORT_148_en = reset;
  assign mem_MPORT_149_data = 20'h0;
  assign mem_MPORT_149_addr = 8'h95;
  assign mem_MPORT_149_mask = 1'h1;
  assign mem_MPORT_149_en = reset;
  assign mem_MPORT_150_data = 20'h0;
  assign mem_MPORT_150_addr = 8'h96;
  assign mem_MPORT_150_mask = 1'h1;
  assign mem_MPORT_150_en = reset;
  assign mem_MPORT_151_data = 20'h0;
  assign mem_MPORT_151_addr = 8'h97;
  assign mem_MPORT_151_mask = 1'h1;
  assign mem_MPORT_151_en = reset;
  assign mem_MPORT_152_data = 20'h0;
  assign mem_MPORT_152_addr = 8'h98;
  assign mem_MPORT_152_mask = 1'h1;
  assign mem_MPORT_152_en = reset;
  assign mem_MPORT_153_data = 20'h0;
  assign mem_MPORT_153_addr = 8'h99;
  assign mem_MPORT_153_mask = 1'h1;
  assign mem_MPORT_153_en = reset;
  assign mem_MPORT_154_data = 20'h0;
  assign mem_MPORT_154_addr = 8'h9a;
  assign mem_MPORT_154_mask = 1'h1;
  assign mem_MPORT_154_en = reset;
  assign mem_MPORT_155_data = 20'h0;
  assign mem_MPORT_155_addr = 8'h9b;
  assign mem_MPORT_155_mask = 1'h1;
  assign mem_MPORT_155_en = reset;
  assign mem_MPORT_156_data = 20'h0;
  assign mem_MPORT_156_addr = 8'h9c;
  assign mem_MPORT_156_mask = 1'h1;
  assign mem_MPORT_156_en = reset;
  assign mem_MPORT_157_data = 20'h0;
  assign mem_MPORT_157_addr = 8'h9d;
  assign mem_MPORT_157_mask = 1'h1;
  assign mem_MPORT_157_en = reset;
  assign mem_MPORT_158_data = 20'h0;
  assign mem_MPORT_158_addr = 8'h9e;
  assign mem_MPORT_158_mask = 1'h1;
  assign mem_MPORT_158_en = reset;
  assign mem_MPORT_159_data = 20'h0;
  assign mem_MPORT_159_addr = 8'h9f;
  assign mem_MPORT_159_mask = 1'h1;
  assign mem_MPORT_159_en = reset;
  assign mem_MPORT_160_data = 20'h0;
  assign mem_MPORT_160_addr = 8'ha0;
  assign mem_MPORT_160_mask = 1'h1;
  assign mem_MPORT_160_en = reset;
  assign mem_MPORT_161_data = 20'h0;
  assign mem_MPORT_161_addr = 8'ha1;
  assign mem_MPORT_161_mask = 1'h1;
  assign mem_MPORT_161_en = reset;
  assign mem_MPORT_162_data = 20'h0;
  assign mem_MPORT_162_addr = 8'ha2;
  assign mem_MPORT_162_mask = 1'h1;
  assign mem_MPORT_162_en = reset;
  assign mem_MPORT_163_data = 20'h0;
  assign mem_MPORT_163_addr = 8'ha3;
  assign mem_MPORT_163_mask = 1'h1;
  assign mem_MPORT_163_en = reset;
  assign mem_MPORT_164_data = 20'h0;
  assign mem_MPORT_164_addr = 8'ha4;
  assign mem_MPORT_164_mask = 1'h1;
  assign mem_MPORT_164_en = reset;
  assign mem_MPORT_165_data = 20'h0;
  assign mem_MPORT_165_addr = 8'ha5;
  assign mem_MPORT_165_mask = 1'h1;
  assign mem_MPORT_165_en = reset;
  assign mem_MPORT_166_data = 20'h0;
  assign mem_MPORT_166_addr = 8'ha6;
  assign mem_MPORT_166_mask = 1'h1;
  assign mem_MPORT_166_en = reset;
  assign mem_MPORT_167_data = 20'h0;
  assign mem_MPORT_167_addr = 8'ha7;
  assign mem_MPORT_167_mask = 1'h1;
  assign mem_MPORT_167_en = reset;
  assign mem_MPORT_168_data = 20'h0;
  assign mem_MPORT_168_addr = 8'ha8;
  assign mem_MPORT_168_mask = 1'h1;
  assign mem_MPORT_168_en = reset;
  assign mem_MPORT_169_data = 20'h0;
  assign mem_MPORT_169_addr = 8'ha9;
  assign mem_MPORT_169_mask = 1'h1;
  assign mem_MPORT_169_en = reset;
  assign mem_MPORT_170_data = 20'h0;
  assign mem_MPORT_170_addr = 8'haa;
  assign mem_MPORT_170_mask = 1'h1;
  assign mem_MPORT_170_en = reset;
  assign mem_MPORT_171_data = 20'h0;
  assign mem_MPORT_171_addr = 8'hab;
  assign mem_MPORT_171_mask = 1'h1;
  assign mem_MPORT_171_en = reset;
  assign mem_MPORT_172_data = 20'h0;
  assign mem_MPORT_172_addr = 8'hac;
  assign mem_MPORT_172_mask = 1'h1;
  assign mem_MPORT_172_en = reset;
  assign mem_MPORT_173_data = 20'h0;
  assign mem_MPORT_173_addr = 8'had;
  assign mem_MPORT_173_mask = 1'h1;
  assign mem_MPORT_173_en = reset;
  assign mem_MPORT_174_data = 20'h0;
  assign mem_MPORT_174_addr = 8'hae;
  assign mem_MPORT_174_mask = 1'h1;
  assign mem_MPORT_174_en = reset;
  assign mem_MPORT_175_data = 20'h0;
  assign mem_MPORT_175_addr = 8'haf;
  assign mem_MPORT_175_mask = 1'h1;
  assign mem_MPORT_175_en = reset;
  assign mem_MPORT_176_data = 20'h0;
  assign mem_MPORT_176_addr = 8'hb0;
  assign mem_MPORT_176_mask = 1'h1;
  assign mem_MPORT_176_en = reset;
  assign mem_MPORT_177_data = 20'h0;
  assign mem_MPORT_177_addr = 8'hb1;
  assign mem_MPORT_177_mask = 1'h1;
  assign mem_MPORT_177_en = reset;
  assign mem_MPORT_178_data = 20'h0;
  assign mem_MPORT_178_addr = 8'hb2;
  assign mem_MPORT_178_mask = 1'h1;
  assign mem_MPORT_178_en = reset;
  assign mem_MPORT_179_data = 20'h0;
  assign mem_MPORT_179_addr = 8'hb3;
  assign mem_MPORT_179_mask = 1'h1;
  assign mem_MPORT_179_en = reset;
  assign mem_MPORT_180_data = 20'h0;
  assign mem_MPORT_180_addr = 8'hb4;
  assign mem_MPORT_180_mask = 1'h1;
  assign mem_MPORT_180_en = reset;
  assign mem_MPORT_181_data = 20'h0;
  assign mem_MPORT_181_addr = 8'hb5;
  assign mem_MPORT_181_mask = 1'h1;
  assign mem_MPORT_181_en = reset;
  assign mem_MPORT_182_data = 20'h0;
  assign mem_MPORT_182_addr = 8'hb6;
  assign mem_MPORT_182_mask = 1'h1;
  assign mem_MPORT_182_en = reset;
  assign mem_MPORT_183_data = 20'h0;
  assign mem_MPORT_183_addr = 8'hb7;
  assign mem_MPORT_183_mask = 1'h1;
  assign mem_MPORT_183_en = reset;
  assign mem_MPORT_184_data = 20'h0;
  assign mem_MPORT_184_addr = 8'hb8;
  assign mem_MPORT_184_mask = 1'h1;
  assign mem_MPORT_184_en = reset;
  assign mem_MPORT_185_data = 20'h0;
  assign mem_MPORT_185_addr = 8'hb9;
  assign mem_MPORT_185_mask = 1'h1;
  assign mem_MPORT_185_en = reset;
  assign mem_MPORT_186_data = 20'h0;
  assign mem_MPORT_186_addr = 8'hba;
  assign mem_MPORT_186_mask = 1'h1;
  assign mem_MPORT_186_en = reset;
  assign mem_MPORT_187_data = 20'h0;
  assign mem_MPORT_187_addr = 8'hbb;
  assign mem_MPORT_187_mask = 1'h1;
  assign mem_MPORT_187_en = reset;
  assign mem_MPORT_188_data = 20'h0;
  assign mem_MPORT_188_addr = 8'hbc;
  assign mem_MPORT_188_mask = 1'h1;
  assign mem_MPORT_188_en = reset;
  assign mem_MPORT_189_data = 20'h0;
  assign mem_MPORT_189_addr = 8'hbd;
  assign mem_MPORT_189_mask = 1'h1;
  assign mem_MPORT_189_en = reset;
  assign mem_MPORT_190_data = 20'h0;
  assign mem_MPORT_190_addr = 8'hbe;
  assign mem_MPORT_190_mask = 1'h1;
  assign mem_MPORT_190_en = reset;
  assign mem_MPORT_191_data = 20'h0;
  assign mem_MPORT_191_addr = 8'hbf;
  assign mem_MPORT_191_mask = 1'h1;
  assign mem_MPORT_191_en = reset;
  assign mem_MPORT_192_data = 20'h0;
  assign mem_MPORT_192_addr = 8'hc0;
  assign mem_MPORT_192_mask = 1'h1;
  assign mem_MPORT_192_en = reset;
  assign mem_MPORT_193_data = 20'h0;
  assign mem_MPORT_193_addr = 8'hc1;
  assign mem_MPORT_193_mask = 1'h1;
  assign mem_MPORT_193_en = reset;
  assign mem_MPORT_194_data = 20'h0;
  assign mem_MPORT_194_addr = 8'hc2;
  assign mem_MPORT_194_mask = 1'h1;
  assign mem_MPORT_194_en = reset;
  assign mem_MPORT_195_data = 20'h0;
  assign mem_MPORT_195_addr = 8'hc3;
  assign mem_MPORT_195_mask = 1'h1;
  assign mem_MPORT_195_en = reset;
  assign mem_MPORT_196_data = 20'h0;
  assign mem_MPORT_196_addr = 8'hc4;
  assign mem_MPORT_196_mask = 1'h1;
  assign mem_MPORT_196_en = reset;
  assign mem_MPORT_197_data = 20'h0;
  assign mem_MPORT_197_addr = 8'hc5;
  assign mem_MPORT_197_mask = 1'h1;
  assign mem_MPORT_197_en = reset;
  assign mem_MPORT_198_data = 20'h0;
  assign mem_MPORT_198_addr = 8'hc6;
  assign mem_MPORT_198_mask = 1'h1;
  assign mem_MPORT_198_en = reset;
  assign mem_MPORT_199_data = 20'h0;
  assign mem_MPORT_199_addr = 8'hc7;
  assign mem_MPORT_199_mask = 1'h1;
  assign mem_MPORT_199_en = reset;
  assign mem_MPORT_200_data = 20'h0;
  assign mem_MPORT_200_addr = 8'hc8;
  assign mem_MPORT_200_mask = 1'h1;
  assign mem_MPORT_200_en = reset;
  assign mem_MPORT_201_data = 20'h0;
  assign mem_MPORT_201_addr = 8'hc9;
  assign mem_MPORT_201_mask = 1'h1;
  assign mem_MPORT_201_en = reset;
  assign mem_MPORT_202_data = 20'h0;
  assign mem_MPORT_202_addr = 8'hca;
  assign mem_MPORT_202_mask = 1'h1;
  assign mem_MPORT_202_en = reset;
  assign mem_MPORT_203_data = 20'h0;
  assign mem_MPORT_203_addr = 8'hcb;
  assign mem_MPORT_203_mask = 1'h1;
  assign mem_MPORT_203_en = reset;
  assign mem_MPORT_204_data = 20'h0;
  assign mem_MPORT_204_addr = 8'hcc;
  assign mem_MPORT_204_mask = 1'h1;
  assign mem_MPORT_204_en = reset;
  assign mem_MPORT_205_data = 20'h0;
  assign mem_MPORT_205_addr = 8'hcd;
  assign mem_MPORT_205_mask = 1'h1;
  assign mem_MPORT_205_en = reset;
  assign mem_MPORT_206_data = 20'h0;
  assign mem_MPORT_206_addr = 8'hce;
  assign mem_MPORT_206_mask = 1'h1;
  assign mem_MPORT_206_en = reset;
  assign mem_MPORT_207_data = 20'h0;
  assign mem_MPORT_207_addr = 8'hcf;
  assign mem_MPORT_207_mask = 1'h1;
  assign mem_MPORT_207_en = reset;
  assign mem_MPORT_208_data = 20'h0;
  assign mem_MPORT_208_addr = 8'hd0;
  assign mem_MPORT_208_mask = 1'h1;
  assign mem_MPORT_208_en = reset;
  assign mem_MPORT_209_data = 20'h0;
  assign mem_MPORT_209_addr = 8'hd1;
  assign mem_MPORT_209_mask = 1'h1;
  assign mem_MPORT_209_en = reset;
  assign mem_MPORT_210_data = 20'h0;
  assign mem_MPORT_210_addr = 8'hd2;
  assign mem_MPORT_210_mask = 1'h1;
  assign mem_MPORT_210_en = reset;
  assign mem_MPORT_211_data = 20'h0;
  assign mem_MPORT_211_addr = 8'hd3;
  assign mem_MPORT_211_mask = 1'h1;
  assign mem_MPORT_211_en = reset;
  assign mem_MPORT_212_data = 20'h0;
  assign mem_MPORT_212_addr = 8'hd4;
  assign mem_MPORT_212_mask = 1'h1;
  assign mem_MPORT_212_en = reset;
  assign mem_MPORT_213_data = 20'h0;
  assign mem_MPORT_213_addr = 8'hd5;
  assign mem_MPORT_213_mask = 1'h1;
  assign mem_MPORT_213_en = reset;
  assign mem_MPORT_214_data = 20'h0;
  assign mem_MPORT_214_addr = 8'hd6;
  assign mem_MPORT_214_mask = 1'h1;
  assign mem_MPORT_214_en = reset;
  assign mem_MPORT_215_data = 20'h0;
  assign mem_MPORT_215_addr = 8'hd7;
  assign mem_MPORT_215_mask = 1'h1;
  assign mem_MPORT_215_en = reset;
  assign mem_MPORT_216_data = 20'h0;
  assign mem_MPORT_216_addr = 8'hd8;
  assign mem_MPORT_216_mask = 1'h1;
  assign mem_MPORT_216_en = reset;
  assign mem_MPORT_217_data = 20'h0;
  assign mem_MPORT_217_addr = 8'hd9;
  assign mem_MPORT_217_mask = 1'h1;
  assign mem_MPORT_217_en = reset;
  assign mem_MPORT_218_data = 20'h0;
  assign mem_MPORT_218_addr = 8'hda;
  assign mem_MPORT_218_mask = 1'h1;
  assign mem_MPORT_218_en = reset;
  assign mem_MPORT_219_data = 20'h0;
  assign mem_MPORT_219_addr = 8'hdb;
  assign mem_MPORT_219_mask = 1'h1;
  assign mem_MPORT_219_en = reset;
  assign mem_MPORT_220_data = 20'h0;
  assign mem_MPORT_220_addr = 8'hdc;
  assign mem_MPORT_220_mask = 1'h1;
  assign mem_MPORT_220_en = reset;
  assign mem_MPORT_221_data = 20'h0;
  assign mem_MPORT_221_addr = 8'hdd;
  assign mem_MPORT_221_mask = 1'h1;
  assign mem_MPORT_221_en = reset;
  assign mem_MPORT_222_data = 20'h0;
  assign mem_MPORT_222_addr = 8'hde;
  assign mem_MPORT_222_mask = 1'h1;
  assign mem_MPORT_222_en = reset;
  assign mem_MPORT_223_data = 20'h0;
  assign mem_MPORT_223_addr = 8'hdf;
  assign mem_MPORT_223_mask = 1'h1;
  assign mem_MPORT_223_en = reset;
  assign mem_MPORT_224_data = 20'h0;
  assign mem_MPORT_224_addr = 8'he0;
  assign mem_MPORT_224_mask = 1'h1;
  assign mem_MPORT_224_en = reset;
  assign mem_MPORT_225_data = 20'h0;
  assign mem_MPORT_225_addr = 8'he1;
  assign mem_MPORT_225_mask = 1'h1;
  assign mem_MPORT_225_en = reset;
  assign mem_MPORT_226_data = 20'h0;
  assign mem_MPORT_226_addr = 8'he2;
  assign mem_MPORT_226_mask = 1'h1;
  assign mem_MPORT_226_en = reset;
  assign mem_MPORT_227_data = 20'h0;
  assign mem_MPORT_227_addr = 8'he3;
  assign mem_MPORT_227_mask = 1'h1;
  assign mem_MPORT_227_en = reset;
  assign mem_MPORT_228_data = 20'h0;
  assign mem_MPORT_228_addr = 8'he4;
  assign mem_MPORT_228_mask = 1'h1;
  assign mem_MPORT_228_en = reset;
  assign mem_MPORT_229_data = 20'h0;
  assign mem_MPORT_229_addr = 8'he5;
  assign mem_MPORT_229_mask = 1'h1;
  assign mem_MPORT_229_en = reset;
  assign mem_MPORT_230_data = 20'h0;
  assign mem_MPORT_230_addr = 8'he6;
  assign mem_MPORT_230_mask = 1'h1;
  assign mem_MPORT_230_en = reset;
  assign mem_MPORT_231_data = 20'h0;
  assign mem_MPORT_231_addr = 8'he7;
  assign mem_MPORT_231_mask = 1'h1;
  assign mem_MPORT_231_en = reset;
  assign mem_MPORT_232_data = 20'h0;
  assign mem_MPORT_232_addr = 8'he8;
  assign mem_MPORT_232_mask = 1'h1;
  assign mem_MPORT_232_en = reset;
  assign mem_MPORT_233_data = 20'h0;
  assign mem_MPORT_233_addr = 8'he9;
  assign mem_MPORT_233_mask = 1'h1;
  assign mem_MPORT_233_en = reset;
  assign mem_MPORT_234_data = 20'h0;
  assign mem_MPORT_234_addr = 8'hea;
  assign mem_MPORT_234_mask = 1'h1;
  assign mem_MPORT_234_en = reset;
  assign mem_MPORT_235_data = 20'h0;
  assign mem_MPORT_235_addr = 8'heb;
  assign mem_MPORT_235_mask = 1'h1;
  assign mem_MPORT_235_en = reset;
  assign mem_MPORT_236_data = 20'h0;
  assign mem_MPORT_236_addr = 8'hec;
  assign mem_MPORT_236_mask = 1'h1;
  assign mem_MPORT_236_en = reset;
  assign mem_MPORT_237_data = 20'h0;
  assign mem_MPORT_237_addr = 8'hed;
  assign mem_MPORT_237_mask = 1'h1;
  assign mem_MPORT_237_en = reset;
  assign mem_MPORT_238_data = 20'h0;
  assign mem_MPORT_238_addr = 8'hee;
  assign mem_MPORT_238_mask = 1'h1;
  assign mem_MPORT_238_en = reset;
  assign mem_MPORT_239_data = 20'h0;
  assign mem_MPORT_239_addr = 8'hef;
  assign mem_MPORT_239_mask = 1'h1;
  assign mem_MPORT_239_en = reset;
  assign mem_MPORT_240_data = 20'h0;
  assign mem_MPORT_240_addr = 8'hf0;
  assign mem_MPORT_240_mask = 1'h1;
  assign mem_MPORT_240_en = reset;
  assign mem_MPORT_241_data = 20'h0;
  assign mem_MPORT_241_addr = 8'hf1;
  assign mem_MPORT_241_mask = 1'h1;
  assign mem_MPORT_241_en = reset;
  assign mem_MPORT_242_data = 20'h0;
  assign mem_MPORT_242_addr = 8'hf2;
  assign mem_MPORT_242_mask = 1'h1;
  assign mem_MPORT_242_en = reset;
  assign mem_MPORT_243_data = 20'h0;
  assign mem_MPORT_243_addr = 8'hf3;
  assign mem_MPORT_243_mask = 1'h1;
  assign mem_MPORT_243_en = reset;
  assign mem_MPORT_244_data = 20'h0;
  assign mem_MPORT_244_addr = 8'hf4;
  assign mem_MPORT_244_mask = 1'h1;
  assign mem_MPORT_244_en = reset;
  assign mem_MPORT_245_data = 20'h0;
  assign mem_MPORT_245_addr = 8'hf5;
  assign mem_MPORT_245_mask = 1'h1;
  assign mem_MPORT_245_en = reset;
  assign mem_MPORT_246_data = 20'h0;
  assign mem_MPORT_246_addr = 8'hf6;
  assign mem_MPORT_246_mask = 1'h1;
  assign mem_MPORT_246_en = reset;
  assign mem_MPORT_247_data = 20'h0;
  assign mem_MPORT_247_addr = 8'hf7;
  assign mem_MPORT_247_mask = 1'h1;
  assign mem_MPORT_247_en = reset;
  assign mem_MPORT_248_data = 20'h0;
  assign mem_MPORT_248_addr = 8'hf8;
  assign mem_MPORT_248_mask = 1'h1;
  assign mem_MPORT_248_en = reset;
  assign mem_MPORT_249_data = 20'h0;
  assign mem_MPORT_249_addr = 8'hf9;
  assign mem_MPORT_249_mask = 1'h1;
  assign mem_MPORT_249_en = reset;
  assign mem_MPORT_250_data = 20'h0;
  assign mem_MPORT_250_addr = 8'hfa;
  assign mem_MPORT_250_mask = 1'h1;
  assign mem_MPORT_250_en = reset;
  assign mem_MPORT_251_data = 20'h0;
  assign mem_MPORT_251_addr = 8'hfb;
  assign mem_MPORT_251_mask = 1'h1;
  assign mem_MPORT_251_en = reset;
  assign mem_MPORT_252_data = 20'h0;
  assign mem_MPORT_252_addr = 8'hfc;
  assign mem_MPORT_252_mask = 1'h1;
  assign mem_MPORT_252_en = reset;
  assign mem_MPORT_253_data = 20'h0;
  assign mem_MPORT_253_addr = 8'hfd;
  assign mem_MPORT_253_mask = 1'h1;
  assign mem_MPORT_253_en = reset;
  assign mem_MPORT_254_data = 20'h0;
  assign mem_MPORT_254_addr = 8'hfe;
  assign mem_MPORT_254_mask = 1'h1;
  assign mem_MPORT_254_en = reset;
  assign mem_MPORT_255_data = 20'h0;
  assign mem_MPORT_255_addr = 8'hff;
  assign mem_MPORT_255_mask = 1'h1;
  assign mem_MPORT_255_en = reset;
  assign mem_MPORT_256_data = io_w_data;
  assign mem_MPORT_256_addr = io_w_addr;
  assign mem_MPORT_256_mask = 1'h1;
  assign mem_MPORT_256_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_129_en & mem_MPORT_129_mask) begin
      mem[mem_MPORT_129_addr] <= mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_130_en & mem_MPORT_130_mask) begin
      mem[mem_MPORT_130_addr] <= mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_131_en & mem_MPORT_131_mask) begin
      mem[mem_MPORT_131_addr] <= mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_132_en & mem_MPORT_132_mask) begin
      mem[mem_MPORT_132_addr] <= mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_133_en & mem_MPORT_133_mask) begin
      mem[mem_MPORT_133_addr] <= mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_134_en & mem_MPORT_134_mask) begin
      mem[mem_MPORT_134_addr] <= mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_135_en & mem_MPORT_135_mask) begin
      mem[mem_MPORT_135_addr] <= mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_136_en & mem_MPORT_136_mask) begin
      mem[mem_MPORT_136_addr] <= mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_137_en & mem_MPORT_137_mask) begin
      mem[mem_MPORT_137_addr] <= mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_138_en & mem_MPORT_138_mask) begin
      mem[mem_MPORT_138_addr] <= mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_139_en & mem_MPORT_139_mask) begin
      mem[mem_MPORT_139_addr] <= mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_140_en & mem_MPORT_140_mask) begin
      mem[mem_MPORT_140_addr] <= mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_141_en & mem_MPORT_141_mask) begin
      mem[mem_MPORT_141_addr] <= mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_142_en & mem_MPORT_142_mask) begin
      mem[mem_MPORT_142_addr] <= mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_143_en & mem_MPORT_143_mask) begin
      mem[mem_MPORT_143_addr] <= mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_144_en & mem_MPORT_144_mask) begin
      mem[mem_MPORT_144_addr] <= mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_145_en & mem_MPORT_145_mask) begin
      mem[mem_MPORT_145_addr] <= mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_146_en & mem_MPORT_146_mask) begin
      mem[mem_MPORT_146_addr] <= mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_147_en & mem_MPORT_147_mask) begin
      mem[mem_MPORT_147_addr] <= mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_148_en & mem_MPORT_148_mask) begin
      mem[mem_MPORT_148_addr] <= mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_149_en & mem_MPORT_149_mask) begin
      mem[mem_MPORT_149_addr] <= mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_150_en & mem_MPORT_150_mask) begin
      mem[mem_MPORT_150_addr] <= mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_151_en & mem_MPORT_151_mask) begin
      mem[mem_MPORT_151_addr] <= mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_152_en & mem_MPORT_152_mask) begin
      mem[mem_MPORT_152_addr] <= mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_153_en & mem_MPORT_153_mask) begin
      mem[mem_MPORT_153_addr] <= mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_154_en & mem_MPORT_154_mask) begin
      mem[mem_MPORT_154_addr] <= mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_155_en & mem_MPORT_155_mask) begin
      mem[mem_MPORT_155_addr] <= mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_156_en & mem_MPORT_156_mask) begin
      mem[mem_MPORT_156_addr] <= mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_157_en & mem_MPORT_157_mask) begin
      mem[mem_MPORT_157_addr] <= mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_158_en & mem_MPORT_158_mask) begin
      mem[mem_MPORT_158_addr] <= mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_159_en & mem_MPORT_159_mask) begin
      mem[mem_MPORT_159_addr] <= mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_160_en & mem_MPORT_160_mask) begin
      mem[mem_MPORT_160_addr] <= mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_161_en & mem_MPORT_161_mask) begin
      mem[mem_MPORT_161_addr] <= mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_162_en & mem_MPORT_162_mask) begin
      mem[mem_MPORT_162_addr] <= mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_163_en & mem_MPORT_163_mask) begin
      mem[mem_MPORT_163_addr] <= mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_164_en & mem_MPORT_164_mask) begin
      mem[mem_MPORT_164_addr] <= mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_165_en & mem_MPORT_165_mask) begin
      mem[mem_MPORT_165_addr] <= mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_166_en & mem_MPORT_166_mask) begin
      mem[mem_MPORT_166_addr] <= mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_167_en & mem_MPORT_167_mask) begin
      mem[mem_MPORT_167_addr] <= mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_168_en & mem_MPORT_168_mask) begin
      mem[mem_MPORT_168_addr] <= mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_169_en & mem_MPORT_169_mask) begin
      mem[mem_MPORT_169_addr] <= mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_170_en & mem_MPORT_170_mask) begin
      mem[mem_MPORT_170_addr] <= mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_171_en & mem_MPORT_171_mask) begin
      mem[mem_MPORT_171_addr] <= mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_172_en & mem_MPORT_172_mask) begin
      mem[mem_MPORT_172_addr] <= mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_173_en & mem_MPORT_173_mask) begin
      mem[mem_MPORT_173_addr] <= mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_174_en & mem_MPORT_174_mask) begin
      mem[mem_MPORT_174_addr] <= mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_175_en & mem_MPORT_175_mask) begin
      mem[mem_MPORT_175_addr] <= mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_176_en & mem_MPORT_176_mask) begin
      mem[mem_MPORT_176_addr] <= mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_177_en & mem_MPORT_177_mask) begin
      mem[mem_MPORT_177_addr] <= mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_178_en & mem_MPORT_178_mask) begin
      mem[mem_MPORT_178_addr] <= mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_179_en & mem_MPORT_179_mask) begin
      mem[mem_MPORT_179_addr] <= mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_180_en & mem_MPORT_180_mask) begin
      mem[mem_MPORT_180_addr] <= mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_181_en & mem_MPORT_181_mask) begin
      mem[mem_MPORT_181_addr] <= mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_182_en & mem_MPORT_182_mask) begin
      mem[mem_MPORT_182_addr] <= mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_183_en & mem_MPORT_183_mask) begin
      mem[mem_MPORT_183_addr] <= mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_184_en & mem_MPORT_184_mask) begin
      mem[mem_MPORT_184_addr] <= mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_185_en & mem_MPORT_185_mask) begin
      mem[mem_MPORT_185_addr] <= mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_186_en & mem_MPORT_186_mask) begin
      mem[mem_MPORT_186_addr] <= mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_187_en & mem_MPORT_187_mask) begin
      mem[mem_MPORT_187_addr] <= mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_188_en & mem_MPORT_188_mask) begin
      mem[mem_MPORT_188_addr] <= mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_189_en & mem_MPORT_189_mask) begin
      mem[mem_MPORT_189_addr] <= mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_190_en & mem_MPORT_190_mask) begin
      mem[mem_MPORT_190_addr] <= mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_191_en & mem_MPORT_191_mask) begin
      mem[mem_MPORT_191_addr] <= mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_192_en & mem_MPORT_192_mask) begin
      mem[mem_MPORT_192_addr] <= mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_193_en & mem_MPORT_193_mask) begin
      mem[mem_MPORT_193_addr] <= mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_194_en & mem_MPORT_194_mask) begin
      mem[mem_MPORT_194_addr] <= mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_195_en & mem_MPORT_195_mask) begin
      mem[mem_MPORT_195_addr] <= mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_196_en & mem_MPORT_196_mask) begin
      mem[mem_MPORT_196_addr] <= mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_197_en & mem_MPORT_197_mask) begin
      mem[mem_MPORT_197_addr] <= mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_198_en & mem_MPORT_198_mask) begin
      mem[mem_MPORT_198_addr] <= mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_199_en & mem_MPORT_199_mask) begin
      mem[mem_MPORT_199_addr] <= mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_200_en & mem_MPORT_200_mask) begin
      mem[mem_MPORT_200_addr] <= mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_201_en & mem_MPORT_201_mask) begin
      mem[mem_MPORT_201_addr] <= mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_202_en & mem_MPORT_202_mask) begin
      mem[mem_MPORT_202_addr] <= mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_203_en & mem_MPORT_203_mask) begin
      mem[mem_MPORT_203_addr] <= mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_204_en & mem_MPORT_204_mask) begin
      mem[mem_MPORT_204_addr] <= mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_205_en & mem_MPORT_205_mask) begin
      mem[mem_MPORT_205_addr] <= mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_206_en & mem_MPORT_206_mask) begin
      mem[mem_MPORT_206_addr] <= mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_207_en & mem_MPORT_207_mask) begin
      mem[mem_MPORT_207_addr] <= mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_208_en & mem_MPORT_208_mask) begin
      mem[mem_MPORT_208_addr] <= mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_209_en & mem_MPORT_209_mask) begin
      mem[mem_MPORT_209_addr] <= mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_210_en & mem_MPORT_210_mask) begin
      mem[mem_MPORT_210_addr] <= mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_211_en & mem_MPORT_211_mask) begin
      mem[mem_MPORT_211_addr] <= mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_212_en & mem_MPORT_212_mask) begin
      mem[mem_MPORT_212_addr] <= mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_213_en & mem_MPORT_213_mask) begin
      mem[mem_MPORT_213_addr] <= mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_214_en & mem_MPORT_214_mask) begin
      mem[mem_MPORT_214_addr] <= mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_215_en & mem_MPORT_215_mask) begin
      mem[mem_MPORT_215_addr] <= mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_216_en & mem_MPORT_216_mask) begin
      mem[mem_MPORT_216_addr] <= mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_217_en & mem_MPORT_217_mask) begin
      mem[mem_MPORT_217_addr] <= mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_218_en & mem_MPORT_218_mask) begin
      mem[mem_MPORT_218_addr] <= mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_219_en & mem_MPORT_219_mask) begin
      mem[mem_MPORT_219_addr] <= mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_220_en & mem_MPORT_220_mask) begin
      mem[mem_MPORT_220_addr] <= mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_221_en & mem_MPORT_221_mask) begin
      mem[mem_MPORT_221_addr] <= mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_222_en & mem_MPORT_222_mask) begin
      mem[mem_MPORT_222_addr] <= mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_223_en & mem_MPORT_223_mask) begin
      mem[mem_MPORT_223_addr] <= mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_224_en & mem_MPORT_224_mask) begin
      mem[mem_MPORT_224_addr] <= mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_225_en & mem_MPORT_225_mask) begin
      mem[mem_MPORT_225_addr] <= mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_226_en & mem_MPORT_226_mask) begin
      mem[mem_MPORT_226_addr] <= mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_227_en & mem_MPORT_227_mask) begin
      mem[mem_MPORT_227_addr] <= mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_228_en & mem_MPORT_228_mask) begin
      mem[mem_MPORT_228_addr] <= mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_229_en & mem_MPORT_229_mask) begin
      mem[mem_MPORT_229_addr] <= mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_230_en & mem_MPORT_230_mask) begin
      mem[mem_MPORT_230_addr] <= mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_231_en & mem_MPORT_231_mask) begin
      mem[mem_MPORT_231_addr] <= mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_232_en & mem_MPORT_232_mask) begin
      mem[mem_MPORT_232_addr] <= mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_233_en & mem_MPORT_233_mask) begin
      mem[mem_MPORT_233_addr] <= mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_234_en & mem_MPORT_234_mask) begin
      mem[mem_MPORT_234_addr] <= mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_235_en & mem_MPORT_235_mask) begin
      mem[mem_MPORT_235_addr] <= mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_236_en & mem_MPORT_236_mask) begin
      mem[mem_MPORT_236_addr] <= mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_237_en & mem_MPORT_237_mask) begin
      mem[mem_MPORT_237_addr] <= mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_238_en & mem_MPORT_238_mask) begin
      mem[mem_MPORT_238_addr] <= mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_239_en & mem_MPORT_239_mask) begin
      mem[mem_MPORT_239_addr] <= mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_240_en & mem_MPORT_240_mask) begin
      mem[mem_MPORT_240_addr] <= mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_241_en & mem_MPORT_241_mask) begin
      mem[mem_MPORT_241_addr] <= mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_242_en & mem_MPORT_242_mask) begin
      mem[mem_MPORT_242_addr] <= mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_243_en & mem_MPORT_243_mask) begin
      mem[mem_MPORT_243_addr] <= mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_244_en & mem_MPORT_244_mask) begin
      mem[mem_MPORT_244_addr] <= mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_245_en & mem_MPORT_245_mask) begin
      mem[mem_MPORT_245_addr] <= mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_246_en & mem_MPORT_246_mask) begin
      mem[mem_MPORT_246_addr] <= mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_247_en & mem_MPORT_247_mask) begin
      mem[mem_MPORT_247_addr] <= mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_248_en & mem_MPORT_248_mask) begin
      mem[mem_MPORT_248_addr] <= mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_249_en & mem_MPORT_249_mask) begin
      mem[mem_MPORT_249_addr] <= mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_250_en & mem_MPORT_250_mask) begin
      mem[mem_MPORT_250_addr] <= mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_251_en & mem_MPORT_251_mask) begin
      mem[mem_MPORT_251_addr] <= mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_252_en & mem_MPORT_252_mask) begin
      mem[mem_MPORT_252_addr] <= mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_253_en & mem_MPORT_253_mask) begin
      mem[mem_MPORT_253_addr] <= mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_254_en & mem_MPORT_254_mask) begin
      mem[mem_MPORT_254_addr] <= mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_255_en & mem_MPORT_255_mask) begin
      mem[mem_MPORT_255_addr] <= mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_256_en & mem_MPORT_256_mask) begin
      mem[mem_MPORT_256_addr] <= mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _RAND_0[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
