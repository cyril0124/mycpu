module BankRam1P_1_53(
  input        clock,
  input        reset,
  input  [7:0] io_addr,
  input        io_rw,
  input  [7:0] io_wdata,
  input  [3:0] io_wmask,
  output [7:0] io_rdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_0 [0:255]; // @[SRAM.scala 36:26]
  wire  ram_0_io_rdata_MPORT_en; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_io_rdata_MPORT_addr; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_io_rdata_MPORT_data; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_1_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_1_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_1_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_1_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_2_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_2_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_2_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_2_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_3_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_3_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_3_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_3_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_4_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_4_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_4_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_4_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_5_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_5_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_5_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_5_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_6_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_6_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_6_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_6_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_7_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_7_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_7_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_7_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_8_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_8_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_8_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_8_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_9_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_9_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_9_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_9_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_10_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_10_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_10_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_10_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_11_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_11_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_11_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_11_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_12_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_12_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_12_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_12_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_13_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_13_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_13_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_13_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_14_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_14_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_14_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_14_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_15_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_15_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_15_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_15_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_16_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_16_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_16_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_16_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_17_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_17_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_17_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_17_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_18_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_18_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_18_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_18_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_19_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_19_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_19_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_19_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_20_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_20_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_20_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_20_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_21_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_21_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_21_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_21_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_22_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_22_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_22_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_22_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_23_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_23_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_23_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_23_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_24_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_24_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_24_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_24_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_25_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_25_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_25_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_25_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_26_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_26_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_26_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_26_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_27_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_27_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_27_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_27_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_28_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_28_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_28_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_28_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_29_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_29_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_29_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_29_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_30_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_30_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_30_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_30_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_31_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_31_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_31_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_31_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_32_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_32_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_32_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_32_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_33_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_33_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_33_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_33_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_34_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_34_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_34_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_34_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_35_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_35_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_35_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_35_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_36_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_36_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_36_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_36_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_37_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_37_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_37_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_37_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_38_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_38_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_38_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_38_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_39_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_39_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_39_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_39_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_40_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_40_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_40_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_40_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_41_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_41_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_41_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_41_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_42_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_42_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_42_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_42_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_43_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_43_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_43_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_43_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_44_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_44_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_44_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_44_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_45_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_45_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_45_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_45_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_46_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_46_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_46_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_46_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_47_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_47_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_47_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_47_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_48_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_48_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_48_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_48_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_49_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_49_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_49_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_49_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_50_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_50_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_50_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_50_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_51_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_51_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_51_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_51_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_52_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_52_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_52_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_52_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_53_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_53_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_53_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_53_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_54_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_54_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_54_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_54_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_55_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_55_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_55_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_55_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_56_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_56_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_56_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_56_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_57_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_57_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_57_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_57_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_58_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_58_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_58_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_58_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_59_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_59_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_59_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_59_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_60_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_60_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_60_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_60_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_61_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_61_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_61_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_61_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_62_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_62_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_62_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_62_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_63_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_63_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_63_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_63_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_64_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_64_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_64_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_64_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_65_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_65_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_65_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_65_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_66_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_66_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_66_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_66_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_67_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_67_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_67_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_67_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_68_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_68_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_68_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_68_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_69_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_69_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_69_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_69_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_70_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_70_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_70_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_70_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_71_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_71_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_71_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_71_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_72_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_72_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_72_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_72_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_73_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_73_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_73_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_73_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_74_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_74_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_74_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_74_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_75_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_75_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_75_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_75_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_76_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_76_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_76_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_76_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_77_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_77_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_77_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_77_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_78_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_78_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_78_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_78_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_79_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_79_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_79_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_79_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_80_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_80_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_80_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_80_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_81_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_81_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_81_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_81_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_82_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_82_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_82_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_82_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_83_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_83_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_83_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_83_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_84_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_84_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_84_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_84_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_85_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_85_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_85_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_85_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_86_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_86_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_86_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_86_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_87_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_87_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_87_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_87_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_88_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_88_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_88_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_88_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_89_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_89_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_89_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_89_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_90_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_90_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_90_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_90_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_91_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_91_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_91_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_91_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_92_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_92_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_92_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_92_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_93_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_93_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_93_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_93_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_94_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_94_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_94_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_94_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_95_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_95_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_95_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_95_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_96_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_96_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_96_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_96_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_97_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_97_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_97_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_97_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_98_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_98_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_98_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_98_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_99_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_99_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_99_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_99_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_100_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_100_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_100_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_100_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_101_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_101_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_101_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_101_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_102_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_102_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_102_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_102_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_103_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_103_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_103_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_103_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_104_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_104_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_104_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_104_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_105_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_105_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_105_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_105_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_106_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_106_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_106_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_106_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_107_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_107_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_107_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_107_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_108_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_108_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_108_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_108_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_109_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_109_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_109_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_109_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_110_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_110_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_110_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_110_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_111_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_111_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_111_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_111_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_112_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_112_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_112_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_112_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_113_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_113_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_113_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_113_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_114_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_114_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_114_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_114_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_115_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_115_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_115_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_115_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_116_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_116_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_116_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_116_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_117_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_117_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_117_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_117_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_118_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_118_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_118_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_118_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_119_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_119_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_119_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_119_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_120_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_120_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_120_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_120_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_121_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_121_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_121_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_121_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_122_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_122_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_122_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_122_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_123_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_123_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_123_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_123_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_124_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_124_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_124_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_124_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_125_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_125_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_125_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_125_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_126_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_126_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_126_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_126_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_127_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_127_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_127_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_127_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_128_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_128_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_128_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_128_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_129_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_129_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_129_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_129_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_130_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_130_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_130_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_130_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_131_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_131_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_131_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_131_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_132_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_132_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_132_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_132_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_133_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_133_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_133_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_133_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_134_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_134_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_134_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_134_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_135_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_135_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_135_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_135_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_136_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_136_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_136_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_136_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_137_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_137_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_137_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_137_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_138_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_138_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_138_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_138_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_139_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_139_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_139_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_139_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_140_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_140_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_140_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_140_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_141_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_141_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_141_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_141_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_142_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_142_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_142_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_142_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_143_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_143_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_143_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_143_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_144_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_144_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_144_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_144_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_145_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_145_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_145_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_145_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_146_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_146_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_146_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_146_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_147_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_147_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_147_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_147_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_148_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_148_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_148_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_148_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_149_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_149_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_149_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_149_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_150_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_150_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_150_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_150_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_151_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_151_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_151_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_151_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_152_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_152_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_152_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_152_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_153_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_153_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_153_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_153_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_154_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_154_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_154_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_154_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_155_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_155_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_155_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_155_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_156_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_156_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_156_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_156_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_157_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_157_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_157_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_157_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_158_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_158_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_158_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_158_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_159_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_159_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_159_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_159_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_160_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_160_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_160_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_160_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_161_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_161_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_161_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_161_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_162_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_162_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_162_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_162_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_163_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_163_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_163_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_163_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_164_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_164_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_164_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_164_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_165_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_165_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_165_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_165_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_166_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_166_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_166_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_166_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_167_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_167_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_167_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_167_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_168_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_168_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_168_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_168_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_169_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_169_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_169_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_169_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_170_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_170_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_170_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_170_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_171_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_171_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_171_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_171_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_172_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_172_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_172_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_172_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_173_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_173_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_173_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_173_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_174_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_174_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_174_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_174_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_175_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_175_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_175_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_175_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_176_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_176_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_176_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_176_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_177_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_177_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_177_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_177_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_178_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_178_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_178_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_178_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_179_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_179_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_179_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_179_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_180_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_180_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_180_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_180_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_181_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_181_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_181_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_181_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_182_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_182_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_182_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_182_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_183_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_183_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_183_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_183_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_184_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_184_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_184_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_184_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_185_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_185_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_185_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_185_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_186_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_186_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_186_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_186_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_187_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_187_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_187_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_187_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_188_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_188_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_188_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_188_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_189_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_189_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_189_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_189_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_190_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_190_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_190_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_190_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_191_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_191_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_191_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_191_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_192_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_192_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_192_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_192_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_193_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_193_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_193_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_193_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_194_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_194_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_194_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_194_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_195_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_195_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_195_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_195_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_196_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_196_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_196_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_196_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_197_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_197_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_197_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_197_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_198_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_198_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_198_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_198_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_199_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_199_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_199_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_199_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_200_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_200_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_200_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_200_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_201_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_201_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_201_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_201_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_202_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_202_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_202_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_202_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_203_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_203_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_203_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_203_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_204_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_204_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_204_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_204_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_205_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_205_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_205_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_205_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_206_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_206_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_206_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_206_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_207_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_207_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_207_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_207_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_208_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_208_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_208_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_208_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_209_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_209_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_209_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_209_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_210_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_210_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_210_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_210_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_211_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_211_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_211_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_211_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_212_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_212_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_212_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_212_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_213_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_213_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_213_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_213_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_214_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_214_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_214_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_214_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_215_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_215_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_215_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_215_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_216_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_216_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_216_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_216_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_217_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_217_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_217_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_217_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_218_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_218_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_218_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_218_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_219_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_219_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_219_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_219_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_220_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_220_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_220_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_220_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_221_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_221_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_221_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_221_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_222_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_222_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_222_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_222_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_223_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_223_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_223_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_223_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_224_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_224_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_224_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_224_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_225_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_225_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_225_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_225_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_226_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_226_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_226_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_226_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_227_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_227_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_227_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_227_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_228_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_228_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_228_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_228_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_229_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_229_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_229_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_229_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_230_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_230_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_230_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_230_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_231_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_231_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_231_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_231_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_232_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_232_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_232_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_232_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_233_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_233_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_233_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_233_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_234_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_234_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_234_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_234_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_235_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_235_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_235_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_235_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_236_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_236_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_236_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_236_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_237_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_237_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_237_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_237_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_238_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_238_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_238_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_238_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_239_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_239_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_239_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_239_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_240_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_240_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_240_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_240_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_241_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_241_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_241_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_241_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_242_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_242_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_242_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_242_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_243_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_243_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_243_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_243_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_244_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_244_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_244_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_244_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_245_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_245_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_245_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_245_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_246_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_246_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_246_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_246_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_247_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_247_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_247_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_247_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_248_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_248_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_248_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_248_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_249_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_249_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_249_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_249_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_250_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_250_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_250_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_250_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_251_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_251_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_251_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_251_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_252_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_252_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_252_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_252_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_253_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_253_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_253_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_253_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_254_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_254_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_254_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_254_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_255_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_255_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_255_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_255_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_0_MPORT_256_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_0_MPORT_256_addr; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_256_mask; // @[SRAM.scala 36:26]
  wire  ram_0_MPORT_256_en; // @[SRAM.scala 36:26]
  reg  ram_0_io_rdata_MPORT_en_pipe_0;
  reg [7:0] ram_0_io_rdata_MPORT_addr_pipe_0;
  reg [1:0] ram_1 [0:255]; // @[SRAM.scala 36:26]
  wire  ram_1_io_rdata_MPORT_en; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_io_rdata_MPORT_addr; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_io_rdata_MPORT_data; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_1_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_1_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_1_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_1_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_2_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_2_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_2_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_2_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_3_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_3_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_3_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_3_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_4_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_4_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_4_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_4_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_5_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_5_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_5_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_5_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_6_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_6_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_6_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_6_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_7_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_7_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_7_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_7_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_8_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_8_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_8_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_8_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_9_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_9_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_9_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_9_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_10_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_10_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_10_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_10_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_11_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_11_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_11_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_11_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_12_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_12_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_12_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_12_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_13_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_13_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_13_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_13_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_14_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_14_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_14_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_14_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_15_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_15_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_15_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_15_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_16_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_16_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_16_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_16_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_17_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_17_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_17_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_17_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_18_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_18_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_18_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_18_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_19_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_19_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_19_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_19_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_20_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_20_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_20_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_20_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_21_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_21_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_21_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_21_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_22_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_22_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_22_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_22_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_23_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_23_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_23_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_23_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_24_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_24_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_24_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_24_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_25_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_25_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_25_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_25_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_26_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_26_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_26_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_26_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_27_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_27_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_27_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_27_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_28_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_28_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_28_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_28_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_29_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_29_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_29_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_29_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_30_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_30_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_30_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_30_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_31_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_31_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_31_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_31_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_32_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_32_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_32_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_32_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_33_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_33_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_33_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_33_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_34_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_34_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_34_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_34_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_35_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_35_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_35_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_35_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_36_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_36_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_36_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_36_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_37_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_37_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_37_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_37_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_38_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_38_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_38_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_38_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_39_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_39_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_39_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_39_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_40_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_40_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_40_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_40_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_41_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_41_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_41_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_41_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_42_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_42_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_42_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_42_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_43_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_43_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_43_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_43_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_44_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_44_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_44_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_44_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_45_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_45_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_45_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_45_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_46_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_46_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_46_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_46_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_47_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_47_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_47_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_47_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_48_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_48_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_48_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_48_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_49_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_49_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_49_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_49_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_50_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_50_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_50_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_50_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_51_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_51_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_51_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_51_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_52_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_52_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_52_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_52_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_53_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_53_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_53_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_53_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_54_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_54_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_54_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_54_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_55_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_55_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_55_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_55_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_56_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_56_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_56_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_56_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_57_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_57_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_57_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_57_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_58_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_58_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_58_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_58_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_59_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_59_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_59_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_59_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_60_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_60_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_60_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_60_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_61_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_61_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_61_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_61_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_62_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_62_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_62_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_62_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_63_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_63_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_63_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_63_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_64_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_64_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_64_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_64_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_65_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_65_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_65_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_65_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_66_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_66_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_66_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_66_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_67_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_67_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_67_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_67_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_68_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_68_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_68_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_68_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_69_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_69_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_69_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_69_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_70_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_70_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_70_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_70_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_71_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_71_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_71_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_71_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_72_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_72_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_72_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_72_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_73_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_73_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_73_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_73_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_74_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_74_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_74_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_74_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_75_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_75_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_75_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_75_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_76_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_76_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_76_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_76_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_77_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_77_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_77_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_77_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_78_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_78_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_78_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_78_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_79_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_79_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_79_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_79_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_80_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_80_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_80_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_80_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_81_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_81_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_81_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_81_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_82_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_82_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_82_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_82_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_83_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_83_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_83_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_83_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_84_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_84_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_84_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_84_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_85_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_85_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_85_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_85_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_86_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_86_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_86_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_86_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_87_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_87_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_87_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_87_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_88_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_88_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_88_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_88_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_89_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_89_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_89_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_89_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_90_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_90_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_90_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_90_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_91_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_91_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_91_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_91_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_92_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_92_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_92_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_92_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_93_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_93_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_93_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_93_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_94_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_94_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_94_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_94_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_95_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_95_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_95_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_95_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_96_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_96_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_96_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_96_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_97_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_97_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_97_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_97_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_98_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_98_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_98_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_98_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_99_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_99_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_99_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_99_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_100_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_100_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_100_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_100_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_101_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_101_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_101_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_101_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_102_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_102_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_102_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_102_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_103_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_103_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_103_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_103_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_104_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_104_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_104_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_104_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_105_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_105_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_105_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_105_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_106_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_106_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_106_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_106_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_107_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_107_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_107_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_107_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_108_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_108_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_108_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_108_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_109_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_109_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_109_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_109_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_110_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_110_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_110_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_110_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_111_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_111_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_111_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_111_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_112_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_112_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_112_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_112_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_113_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_113_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_113_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_113_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_114_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_114_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_114_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_114_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_115_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_115_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_115_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_115_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_116_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_116_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_116_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_116_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_117_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_117_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_117_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_117_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_118_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_118_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_118_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_118_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_119_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_119_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_119_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_119_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_120_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_120_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_120_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_120_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_121_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_121_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_121_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_121_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_122_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_122_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_122_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_122_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_123_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_123_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_123_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_123_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_124_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_124_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_124_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_124_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_125_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_125_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_125_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_125_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_126_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_126_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_126_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_126_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_127_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_127_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_127_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_127_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_128_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_128_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_128_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_128_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_129_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_129_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_129_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_129_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_130_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_130_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_130_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_130_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_131_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_131_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_131_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_131_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_132_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_132_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_132_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_132_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_133_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_133_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_133_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_133_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_134_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_134_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_134_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_134_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_135_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_135_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_135_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_135_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_136_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_136_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_136_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_136_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_137_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_137_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_137_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_137_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_138_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_138_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_138_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_138_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_139_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_139_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_139_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_139_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_140_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_140_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_140_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_140_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_141_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_141_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_141_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_141_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_142_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_142_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_142_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_142_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_143_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_143_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_143_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_143_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_144_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_144_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_144_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_144_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_145_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_145_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_145_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_145_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_146_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_146_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_146_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_146_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_147_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_147_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_147_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_147_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_148_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_148_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_148_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_148_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_149_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_149_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_149_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_149_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_150_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_150_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_150_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_150_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_151_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_151_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_151_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_151_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_152_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_152_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_152_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_152_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_153_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_153_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_153_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_153_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_154_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_154_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_154_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_154_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_155_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_155_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_155_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_155_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_156_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_156_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_156_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_156_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_157_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_157_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_157_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_157_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_158_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_158_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_158_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_158_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_159_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_159_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_159_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_159_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_160_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_160_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_160_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_160_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_161_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_161_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_161_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_161_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_162_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_162_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_162_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_162_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_163_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_163_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_163_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_163_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_164_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_164_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_164_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_164_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_165_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_165_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_165_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_165_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_166_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_166_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_166_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_166_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_167_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_167_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_167_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_167_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_168_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_168_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_168_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_168_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_169_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_169_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_169_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_169_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_170_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_170_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_170_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_170_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_171_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_171_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_171_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_171_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_172_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_172_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_172_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_172_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_173_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_173_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_173_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_173_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_174_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_174_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_174_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_174_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_175_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_175_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_175_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_175_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_176_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_176_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_176_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_176_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_177_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_177_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_177_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_177_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_178_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_178_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_178_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_178_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_179_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_179_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_179_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_179_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_180_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_180_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_180_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_180_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_181_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_181_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_181_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_181_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_182_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_182_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_182_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_182_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_183_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_183_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_183_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_183_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_184_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_184_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_184_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_184_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_185_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_185_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_185_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_185_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_186_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_186_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_186_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_186_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_187_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_187_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_187_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_187_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_188_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_188_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_188_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_188_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_189_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_189_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_189_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_189_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_190_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_190_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_190_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_190_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_191_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_191_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_191_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_191_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_192_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_192_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_192_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_192_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_193_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_193_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_193_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_193_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_194_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_194_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_194_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_194_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_195_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_195_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_195_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_195_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_196_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_196_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_196_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_196_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_197_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_197_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_197_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_197_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_198_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_198_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_198_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_198_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_199_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_199_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_199_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_199_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_200_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_200_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_200_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_200_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_201_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_201_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_201_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_201_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_202_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_202_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_202_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_202_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_203_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_203_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_203_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_203_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_204_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_204_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_204_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_204_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_205_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_205_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_205_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_205_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_206_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_206_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_206_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_206_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_207_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_207_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_207_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_207_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_208_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_208_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_208_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_208_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_209_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_209_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_209_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_209_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_210_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_210_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_210_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_210_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_211_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_211_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_211_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_211_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_212_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_212_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_212_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_212_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_213_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_213_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_213_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_213_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_214_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_214_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_214_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_214_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_215_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_215_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_215_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_215_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_216_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_216_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_216_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_216_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_217_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_217_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_217_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_217_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_218_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_218_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_218_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_218_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_219_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_219_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_219_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_219_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_220_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_220_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_220_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_220_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_221_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_221_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_221_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_221_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_222_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_222_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_222_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_222_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_223_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_223_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_223_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_223_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_224_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_224_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_224_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_224_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_225_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_225_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_225_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_225_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_226_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_226_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_226_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_226_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_227_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_227_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_227_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_227_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_228_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_228_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_228_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_228_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_229_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_229_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_229_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_229_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_230_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_230_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_230_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_230_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_231_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_231_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_231_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_231_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_232_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_232_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_232_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_232_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_233_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_233_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_233_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_233_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_234_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_234_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_234_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_234_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_235_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_235_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_235_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_235_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_236_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_236_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_236_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_236_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_237_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_237_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_237_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_237_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_238_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_238_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_238_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_238_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_239_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_239_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_239_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_239_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_240_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_240_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_240_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_240_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_241_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_241_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_241_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_241_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_242_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_242_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_242_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_242_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_243_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_243_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_243_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_243_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_244_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_244_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_244_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_244_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_245_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_245_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_245_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_245_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_246_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_246_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_246_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_246_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_247_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_247_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_247_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_247_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_248_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_248_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_248_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_248_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_249_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_249_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_249_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_249_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_250_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_250_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_250_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_250_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_251_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_251_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_251_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_251_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_252_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_252_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_252_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_252_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_253_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_253_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_253_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_253_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_254_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_254_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_254_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_254_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_255_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_255_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_255_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_255_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_1_MPORT_256_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_1_MPORT_256_addr; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_256_mask; // @[SRAM.scala 36:26]
  wire  ram_1_MPORT_256_en; // @[SRAM.scala 36:26]
  reg  ram_1_io_rdata_MPORT_en_pipe_0;
  reg [7:0] ram_1_io_rdata_MPORT_addr_pipe_0;
  reg [1:0] ram_2 [0:255]; // @[SRAM.scala 36:26]
  wire  ram_2_io_rdata_MPORT_en; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_io_rdata_MPORT_addr; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_io_rdata_MPORT_data; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_1_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_1_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_1_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_1_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_2_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_2_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_2_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_2_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_3_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_3_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_3_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_3_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_4_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_4_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_4_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_4_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_5_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_5_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_5_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_5_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_6_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_6_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_6_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_6_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_7_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_7_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_7_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_7_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_8_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_8_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_8_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_8_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_9_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_9_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_9_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_9_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_10_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_10_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_10_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_10_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_11_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_11_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_11_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_11_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_12_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_12_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_12_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_12_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_13_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_13_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_13_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_13_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_14_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_14_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_14_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_14_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_15_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_15_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_15_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_15_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_16_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_16_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_16_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_16_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_17_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_17_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_17_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_17_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_18_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_18_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_18_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_18_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_19_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_19_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_19_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_19_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_20_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_20_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_20_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_20_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_21_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_21_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_21_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_21_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_22_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_22_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_22_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_22_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_23_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_23_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_23_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_23_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_24_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_24_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_24_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_24_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_25_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_25_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_25_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_25_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_26_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_26_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_26_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_26_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_27_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_27_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_27_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_27_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_28_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_28_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_28_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_28_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_29_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_29_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_29_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_29_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_30_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_30_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_30_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_30_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_31_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_31_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_31_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_31_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_32_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_32_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_32_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_32_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_33_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_33_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_33_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_33_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_34_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_34_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_34_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_34_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_35_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_35_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_35_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_35_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_36_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_36_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_36_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_36_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_37_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_37_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_37_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_37_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_38_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_38_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_38_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_38_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_39_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_39_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_39_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_39_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_40_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_40_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_40_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_40_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_41_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_41_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_41_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_41_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_42_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_42_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_42_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_42_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_43_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_43_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_43_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_43_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_44_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_44_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_44_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_44_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_45_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_45_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_45_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_45_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_46_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_46_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_46_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_46_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_47_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_47_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_47_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_47_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_48_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_48_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_48_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_48_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_49_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_49_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_49_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_49_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_50_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_50_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_50_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_50_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_51_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_51_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_51_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_51_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_52_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_52_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_52_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_52_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_53_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_53_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_53_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_53_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_54_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_54_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_54_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_54_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_55_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_55_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_55_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_55_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_56_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_56_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_56_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_56_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_57_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_57_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_57_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_57_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_58_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_58_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_58_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_58_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_59_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_59_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_59_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_59_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_60_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_60_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_60_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_60_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_61_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_61_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_61_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_61_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_62_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_62_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_62_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_62_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_63_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_63_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_63_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_63_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_64_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_64_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_64_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_64_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_65_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_65_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_65_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_65_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_66_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_66_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_66_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_66_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_67_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_67_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_67_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_67_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_68_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_68_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_68_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_68_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_69_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_69_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_69_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_69_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_70_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_70_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_70_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_70_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_71_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_71_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_71_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_71_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_72_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_72_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_72_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_72_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_73_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_73_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_73_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_73_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_74_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_74_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_74_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_74_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_75_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_75_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_75_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_75_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_76_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_76_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_76_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_76_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_77_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_77_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_77_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_77_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_78_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_78_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_78_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_78_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_79_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_79_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_79_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_79_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_80_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_80_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_80_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_80_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_81_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_81_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_81_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_81_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_82_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_82_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_82_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_82_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_83_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_83_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_83_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_83_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_84_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_84_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_84_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_84_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_85_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_85_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_85_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_85_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_86_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_86_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_86_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_86_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_87_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_87_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_87_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_87_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_88_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_88_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_88_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_88_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_89_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_89_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_89_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_89_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_90_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_90_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_90_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_90_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_91_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_91_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_91_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_91_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_92_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_92_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_92_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_92_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_93_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_93_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_93_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_93_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_94_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_94_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_94_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_94_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_95_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_95_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_95_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_95_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_96_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_96_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_96_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_96_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_97_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_97_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_97_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_97_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_98_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_98_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_98_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_98_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_99_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_99_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_99_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_99_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_100_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_100_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_100_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_100_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_101_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_101_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_101_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_101_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_102_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_102_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_102_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_102_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_103_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_103_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_103_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_103_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_104_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_104_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_104_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_104_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_105_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_105_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_105_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_105_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_106_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_106_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_106_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_106_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_107_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_107_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_107_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_107_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_108_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_108_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_108_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_108_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_109_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_109_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_109_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_109_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_110_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_110_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_110_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_110_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_111_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_111_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_111_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_111_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_112_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_112_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_112_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_112_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_113_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_113_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_113_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_113_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_114_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_114_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_114_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_114_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_115_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_115_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_115_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_115_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_116_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_116_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_116_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_116_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_117_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_117_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_117_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_117_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_118_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_118_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_118_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_118_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_119_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_119_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_119_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_119_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_120_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_120_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_120_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_120_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_121_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_121_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_121_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_121_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_122_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_122_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_122_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_122_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_123_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_123_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_123_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_123_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_124_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_124_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_124_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_124_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_125_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_125_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_125_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_125_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_126_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_126_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_126_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_126_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_127_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_127_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_127_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_127_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_128_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_128_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_128_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_128_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_129_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_129_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_129_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_129_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_130_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_130_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_130_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_130_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_131_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_131_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_131_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_131_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_132_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_132_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_132_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_132_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_133_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_133_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_133_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_133_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_134_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_134_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_134_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_134_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_135_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_135_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_135_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_135_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_136_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_136_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_136_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_136_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_137_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_137_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_137_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_137_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_138_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_138_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_138_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_138_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_139_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_139_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_139_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_139_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_140_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_140_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_140_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_140_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_141_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_141_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_141_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_141_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_142_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_142_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_142_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_142_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_143_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_143_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_143_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_143_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_144_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_144_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_144_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_144_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_145_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_145_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_145_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_145_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_146_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_146_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_146_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_146_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_147_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_147_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_147_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_147_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_148_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_148_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_148_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_148_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_149_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_149_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_149_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_149_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_150_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_150_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_150_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_150_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_151_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_151_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_151_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_151_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_152_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_152_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_152_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_152_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_153_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_153_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_153_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_153_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_154_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_154_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_154_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_154_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_155_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_155_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_155_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_155_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_156_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_156_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_156_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_156_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_157_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_157_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_157_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_157_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_158_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_158_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_158_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_158_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_159_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_159_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_159_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_159_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_160_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_160_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_160_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_160_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_161_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_161_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_161_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_161_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_162_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_162_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_162_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_162_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_163_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_163_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_163_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_163_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_164_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_164_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_164_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_164_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_165_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_165_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_165_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_165_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_166_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_166_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_166_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_166_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_167_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_167_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_167_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_167_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_168_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_168_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_168_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_168_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_169_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_169_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_169_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_169_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_170_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_170_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_170_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_170_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_171_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_171_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_171_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_171_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_172_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_172_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_172_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_172_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_173_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_173_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_173_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_173_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_174_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_174_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_174_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_174_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_175_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_175_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_175_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_175_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_176_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_176_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_176_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_176_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_177_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_177_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_177_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_177_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_178_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_178_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_178_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_178_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_179_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_179_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_179_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_179_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_180_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_180_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_180_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_180_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_181_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_181_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_181_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_181_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_182_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_182_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_182_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_182_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_183_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_183_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_183_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_183_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_184_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_184_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_184_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_184_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_185_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_185_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_185_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_185_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_186_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_186_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_186_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_186_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_187_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_187_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_187_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_187_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_188_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_188_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_188_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_188_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_189_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_189_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_189_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_189_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_190_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_190_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_190_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_190_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_191_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_191_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_191_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_191_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_192_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_192_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_192_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_192_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_193_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_193_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_193_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_193_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_194_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_194_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_194_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_194_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_195_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_195_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_195_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_195_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_196_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_196_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_196_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_196_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_197_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_197_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_197_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_197_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_198_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_198_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_198_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_198_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_199_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_199_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_199_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_199_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_200_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_200_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_200_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_200_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_201_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_201_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_201_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_201_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_202_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_202_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_202_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_202_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_203_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_203_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_203_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_203_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_204_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_204_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_204_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_204_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_205_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_205_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_205_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_205_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_206_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_206_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_206_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_206_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_207_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_207_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_207_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_207_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_208_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_208_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_208_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_208_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_209_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_209_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_209_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_209_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_210_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_210_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_210_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_210_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_211_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_211_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_211_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_211_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_212_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_212_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_212_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_212_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_213_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_213_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_213_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_213_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_214_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_214_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_214_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_214_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_215_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_215_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_215_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_215_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_216_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_216_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_216_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_216_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_217_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_217_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_217_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_217_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_218_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_218_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_218_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_218_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_219_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_219_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_219_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_219_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_220_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_220_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_220_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_220_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_221_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_221_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_221_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_221_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_222_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_222_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_222_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_222_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_223_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_223_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_223_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_223_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_224_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_224_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_224_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_224_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_225_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_225_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_225_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_225_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_226_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_226_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_226_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_226_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_227_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_227_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_227_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_227_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_228_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_228_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_228_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_228_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_229_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_229_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_229_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_229_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_230_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_230_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_230_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_230_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_231_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_231_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_231_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_231_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_232_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_232_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_232_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_232_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_233_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_233_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_233_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_233_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_234_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_234_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_234_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_234_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_235_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_235_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_235_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_235_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_236_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_236_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_236_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_236_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_237_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_237_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_237_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_237_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_238_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_238_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_238_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_238_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_239_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_239_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_239_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_239_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_240_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_240_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_240_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_240_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_241_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_241_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_241_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_241_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_242_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_242_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_242_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_242_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_243_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_243_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_243_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_243_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_244_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_244_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_244_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_244_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_245_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_245_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_245_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_245_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_246_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_246_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_246_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_246_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_247_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_247_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_247_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_247_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_248_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_248_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_248_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_248_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_249_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_249_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_249_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_249_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_250_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_250_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_250_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_250_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_251_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_251_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_251_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_251_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_252_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_252_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_252_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_252_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_253_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_253_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_253_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_253_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_254_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_254_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_254_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_254_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_255_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_255_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_255_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_255_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_2_MPORT_256_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_2_MPORT_256_addr; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_256_mask; // @[SRAM.scala 36:26]
  wire  ram_2_MPORT_256_en; // @[SRAM.scala 36:26]
  reg  ram_2_io_rdata_MPORT_en_pipe_0;
  reg [7:0] ram_2_io_rdata_MPORT_addr_pipe_0;
  reg [1:0] ram_3 [0:255]; // @[SRAM.scala 36:26]
  wire  ram_3_io_rdata_MPORT_en; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_io_rdata_MPORT_addr; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_io_rdata_MPORT_data; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_1_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_1_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_1_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_1_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_2_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_2_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_2_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_2_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_3_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_3_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_3_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_3_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_4_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_4_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_4_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_4_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_5_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_5_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_5_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_5_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_6_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_6_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_6_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_6_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_7_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_7_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_7_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_7_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_8_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_8_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_8_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_8_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_9_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_9_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_9_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_9_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_10_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_10_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_10_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_10_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_11_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_11_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_11_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_11_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_12_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_12_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_12_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_12_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_13_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_13_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_13_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_13_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_14_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_14_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_14_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_14_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_15_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_15_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_15_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_15_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_16_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_16_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_16_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_16_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_17_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_17_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_17_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_17_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_18_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_18_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_18_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_18_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_19_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_19_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_19_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_19_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_20_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_20_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_20_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_20_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_21_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_21_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_21_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_21_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_22_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_22_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_22_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_22_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_23_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_23_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_23_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_23_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_24_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_24_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_24_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_24_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_25_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_25_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_25_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_25_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_26_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_26_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_26_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_26_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_27_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_27_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_27_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_27_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_28_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_28_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_28_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_28_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_29_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_29_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_29_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_29_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_30_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_30_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_30_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_30_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_31_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_31_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_31_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_31_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_32_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_32_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_32_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_32_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_33_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_33_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_33_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_33_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_34_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_34_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_34_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_34_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_35_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_35_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_35_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_35_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_36_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_36_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_36_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_36_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_37_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_37_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_37_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_37_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_38_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_38_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_38_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_38_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_39_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_39_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_39_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_39_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_40_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_40_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_40_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_40_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_41_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_41_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_41_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_41_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_42_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_42_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_42_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_42_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_43_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_43_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_43_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_43_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_44_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_44_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_44_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_44_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_45_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_45_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_45_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_45_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_46_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_46_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_46_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_46_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_47_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_47_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_47_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_47_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_48_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_48_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_48_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_48_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_49_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_49_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_49_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_49_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_50_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_50_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_50_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_50_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_51_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_51_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_51_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_51_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_52_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_52_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_52_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_52_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_53_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_53_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_53_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_53_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_54_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_54_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_54_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_54_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_55_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_55_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_55_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_55_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_56_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_56_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_56_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_56_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_57_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_57_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_57_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_57_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_58_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_58_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_58_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_58_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_59_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_59_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_59_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_59_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_60_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_60_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_60_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_60_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_61_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_61_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_61_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_61_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_62_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_62_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_62_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_62_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_63_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_63_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_63_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_63_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_64_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_64_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_64_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_64_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_65_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_65_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_65_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_65_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_66_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_66_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_66_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_66_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_67_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_67_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_67_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_67_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_68_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_68_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_68_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_68_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_69_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_69_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_69_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_69_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_70_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_70_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_70_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_70_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_71_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_71_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_71_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_71_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_72_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_72_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_72_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_72_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_73_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_73_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_73_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_73_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_74_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_74_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_74_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_74_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_75_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_75_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_75_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_75_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_76_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_76_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_76_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_76_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_77_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_77_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_77_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_77_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_78_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_78_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_78_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_78_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_79_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_79_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_79_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_79_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_80_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_80_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_80_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_80_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_81_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_81_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_81_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_81_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_82_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_82_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_82_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_82_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_83_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_83_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_83_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_83_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_84_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_84_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_84_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_84_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_85_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_85_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_85_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_85_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_86_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_86_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_86_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_86_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_87_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_87_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_87_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_87_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_88_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_88_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_88_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_88_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_89_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_89_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_89_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_89_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_90_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_90_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_90_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_90_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_91_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_91_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_91_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_91_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_92_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_92_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_92_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_92_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_93_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_93_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_93_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_93_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_94_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_94_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_94_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_94_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_95_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_95_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_95_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_95_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_96_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_96_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_96_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_96_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_97_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_97_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_97_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_97_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_98_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_98_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_98_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_98_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_99_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_99_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_99_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_99_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_100_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_100_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_100_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_100_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_101_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_101_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_101_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_101_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_102_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_102_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_102_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_102_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_103_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_103_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_103_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_103_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_104_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_104_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_104_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_104_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_105_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_105_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_105_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_105_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_106_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_106_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_106_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_106_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_107_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_107_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_107_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_107_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_108_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_108_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_108_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_108_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_109_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_109_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_109_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_109_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_110_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_110_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_110_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_110_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_111_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_111_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_111_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_111_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_112_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_112_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_112_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_112_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_113_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_113_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_113_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_113_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_114_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_114_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_114_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_114_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_115_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_115_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_115_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_115_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_116_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_116_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_116_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_116_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_117_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_117_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_117_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_117_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_118_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_118_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_118_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_118_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_119_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_119_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_119_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_119_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_120_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_120_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_120_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_120_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_121_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_121_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_121_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_121_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_122_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_122_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_122_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_122_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_123_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_123_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_123_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_123_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_124_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_124_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_124_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_124_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_125_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_125_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_125_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_125_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_126_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_126_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_126_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_126_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_127_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_127_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_127_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_127_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_128_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_128_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_128_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_128_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_129_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_129_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_129_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_129_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_130_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_130_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_130_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_130_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_131_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_131_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_131_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_131_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_132_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_132_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_132_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_132_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_133_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_133_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_133_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_133_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_134_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_134_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_134_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_134_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_135_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_135_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_135_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_135_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_136_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_136_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_136_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_136_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_137_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_137_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_137_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_137_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_138_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_138_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_138_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_138_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_139_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_139_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_139_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_139_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_140_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_140_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_140_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_140_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_141_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_141_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_141_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_141_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_142_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_142_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_142_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_142_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_143_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_143_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_143_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_143_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_144_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_144_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_144_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_144_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_145_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_145_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_145_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_145_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_146_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_146_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_146_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_146_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_147_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_147_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_147_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_147_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_148_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_148_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_148_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_148_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_149_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_149_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_149_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_149_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_150_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_150_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_150_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_150_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_151_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_151_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_151_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_151_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_152_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_152_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_152_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_152_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_153_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_153_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_153_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_153_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_154_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_154_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_154_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_154_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_155_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_155_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_155_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_155_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_156_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_156_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_156_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_156_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_157_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_157_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_157_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_157_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_158_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_158_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_158_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_158_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_159_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_159_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_159_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_159_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_160_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_160_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_160_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_160_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_161_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_161_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_161_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_161_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_162_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_162_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_162_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_162_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_163_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_163_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_163_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_163_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_164_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_164_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_164_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_164_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_165_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_165_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_165_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_165_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_166_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_166_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_166_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_166_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_167_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_167_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_167_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_167_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_168_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_168_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_168_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_168_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_169_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_169_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_169_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_169_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_170_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_170_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_170_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_170_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_171_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_171_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_171_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_171_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_172_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_172_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_172_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_172_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_173_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_173_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_173_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_173_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_174_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_174_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_174_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_174_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_175_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_175_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_175_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_175_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_176_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_176_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_176_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_176_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_177_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_177_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_177_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_177_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_178_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_178_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_178_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_178_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_179_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_179_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_179_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_179_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_180_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_180_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_180_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_180_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_181_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_181_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_181_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_181_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_182_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_182_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_182_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_182_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_183_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_183_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_183_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_183_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_184_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_184_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_184_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_184_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_185_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_185_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_185_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_185_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_186_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_186_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_186_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_186_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_187_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_187_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_187_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_187_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_188_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_188_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_188_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_188_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_189_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_189_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_189_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_189_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_190_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_190_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_190_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_190_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_191_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_191_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_191_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_191_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_192_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_192_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_192_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_192_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_193_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_193_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_193_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_193_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_194_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_194_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_194_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_194_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_195_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_195_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_195_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_195_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_196_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_196_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_196_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_196_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_197_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_197_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_197_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_197_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_198_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_198_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_198_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_198_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_199_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_199_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_199_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_199_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_200_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_200_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_200_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_200_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_201_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_201_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_201_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_201_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_202_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_202_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_202_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_202_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_203_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_203_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_203_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_203_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_204_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_204_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_204_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_204_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_205_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_205_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_205_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_205_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_206_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_206_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_206_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_206_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_207_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_207_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_207_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_207_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_208_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_208_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_208_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_208_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_209_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_209_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_209_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_209_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_210_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_210_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_210_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_210_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_211_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_211_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_211_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_211_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_212_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_212_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_212_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_212_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_213_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_213_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_213_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_213_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_214_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_214_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_214_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_214_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_215_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_215_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_215_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_215_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_216_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_216_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_216_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_216_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_217_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_217_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_217_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_217_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_218_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_218_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_218_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_218_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_219_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_219_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_219_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_219_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_220_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_220_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_220_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_220_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_221_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_221_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_221_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_221_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_222_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_222_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_222_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_222_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_223_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_223_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_223_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_223_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_224_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_224_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_224_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_224_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_225_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_225_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_225_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_225_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_226_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_226_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_226_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_226_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_227_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_227_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_227_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_227_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_228_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_228_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_228_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_228_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_229_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_229_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_229_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_229_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_230_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_230_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_230_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_230_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_231_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_231_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_231_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_231_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_232_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_232_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_232_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_232_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_233_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_233_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_233_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_233_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_234_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_234_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_234_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_234_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_235_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_235_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_235_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_235_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_236_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_236_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_236_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_236_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_237_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_237_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_237_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_237_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_238_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_238_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_238_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_238_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_239_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_239_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_239_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_239_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_240_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_240_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_240_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_240_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_241_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_241_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_241_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_241_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_242_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_242_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_242_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_242_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_243_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_243_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_243_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_243_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_244_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_244_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_244_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_244_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_245_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_245_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_245_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_245_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_246_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_246_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_246_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_246_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_247_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_247_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_247_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_247_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_248_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_248_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_248_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_248_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_249_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_249_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_249_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_249_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_250_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_250_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_250_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_250_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_251_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_251_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_251_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_251_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_252_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_252_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_252_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_252_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_253_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_253_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_253_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_253_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_254_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_254_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_254_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_254_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_255_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_255_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_255_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_255_en; // @[SRAM.scala 36:26]
  wire [1:0] ram_3_MPORT_256_data; // @[SRAM.scala 36:26]
  wire [7:0] ram_3_MPORT_256_addr; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_256_mask; // @[SRAM.scala 36:26]
  wire  ram_3_MPORT_256_en; // @[SRAM.scala 36:26]
  reg  ram_3_io_rdata_MPORT_en_pipe_0;
  reg [7:0] ram_3_io_rdata_MPORT_addr_pipe_0;
  wire [3:0] io_rdata_lo = {ram_1_io_rdata_MPORT_data,ram_0_io_rdata_MPORT_data}; // @[SRAM.scala 75:39]
  wire [3:0] io_rdata_hi = {ram_3_io_rdata_MPORT_data,ram_2_io_rdata_MPORT_data}; // @[SRAM.scala 75:39]
  assign ram_0_io_rdata_MPORT_en = ram_0_io_rdata_MPORT_en_pipe_0;
  assign ram_0_io_rdata_MPORT_addr = ram_0_io_rdata_MPORT_addr_pipe_0;
  assign ram_0_io_rdata_MPORT_data = ram_0[ram_0_io_rdata_MPORT_addr]; // @[SRAM.scala 36:26]
  assign ram_0_MPORT_data = 2'h0;
  assign ram_0_MPORT_addr = 8'h0;
  assign ram_0_MPORT_mask = 1'h1;
  assign ram_0_MPORT_en = reset;
  assign ram_0_MPORT_1_data = 2'h0;
  assign ram_0_MPORT_1_addr = 8'h1;
  assign ram_0_MPORT_1_mask = 1'h1;
  assign ram_0_MPORT_1_en = reset;
  assign ram_0_MPORT_2_data = 2'h0;
  assign ram_0_MPORT_2_addr = 8'h2;
  assign ram_0_MPORT_2_mask = 1'h1;
  assign ram_0_MPORT_2_en = reset;
  assign ram_0_MPORT_3_data = 2'h0;
  assign ram_0_MPORT_3_addr = 8'h3;
  assign ram_0_MPORT_3_mask = 1'h1;
  assign ram_0_MPORT_3_en = reset;
  assign ram_0_MPORT_4_data = 2'h0;
  assign ram_0_MPORT_4_addr = 8'h4;
  assign ram_0_MPORT_4_mask = 1'h1;
  assign ram_0_MPORT_4_en = reset;
  assign ram_0_MPORT_5_data = 2'h0;
  assign ram_0_MPORT_5_addr = 8'h5;
  assign ram_0_MPORT_5_mask = 1'h1;
  assign ram_0_MPORT_5_en = reset;
  assign ram_0_MPORT_6_data = 2'h0;
  assign ram_0_MPORT_6_addr = 8'h6;
  assign ram_0_MPORT_6_mask = 1'h1;
  assign ram_0_MPORT_6_en = reset;
  assign ram_0_MPORT_7_data = 2'h0;
  assign ram_0_MPORT_7_addr = 8'h7;
  assign ram_0_MPORT_7_mask = 1'h1;
  assign ram_0_MPORT_7_en = reset;
  assign ram_0_MPORT_8_data = 2'h0;
  assign ram_0_MPORT_8_addr = 8'h8;
  assign ram_0_MPORT_8_mask = 1'h1;
  assign ram_0_MPORT_8_en = reset;
  assign ram_0_MPORT_9_data = 2'h0;
  assign ram_0_MPORT_9_addr = 8'h9;
  assign ram_0_MPORT_9_mask = 1'h1;
  assign ram_0_MPORT_9_en = reset;
  assign ram_0_MPORT_10_data = 2'h0;
  assign ram_0_MPORT_10_addr = 8'ha;
  assign ram_0_MPORT_10_mask = 1'h1;
  assign ram_0_MPORT_10_en = reset;
  assign ram_0_MPORT_11_data = 2'h0;
  assign ram_0_MPORT_11_addr = 8'hb;
  assign ram_0_MPORT_11_mask = 1'h1;
  assign ram_0_MPORT_11_en = reset;
  assign ram_0_MPORT_12_data = 2'h0;
  assign ram_0_MPORT_12_addr = 8'hc;
  assign ram_0_MPORT_12_mask = 1'h1;
  assign ram_0_MPORT_12_en = reset;
  assign ram_0_MPORT_13_data = 2'h0;
  assign ram_0_MPORT_13_addr = 8'hd;
  assign ram_0_MPORT_13_mask = 1'h1;
  assign ram_0_MPORT_13_en = reset;
  assign ram_0_MPORT_14_data = 2'h0;
  assign ram_0_MPORT_14_addr = 8'he;
  assign ram_0_MPORT_14_mask = 1'h1;
  assign ram_0_MPORT_14_en = reset;
  assign ram_0_MPORT_15_data = 2'h0;
  assign ram_0_MPORT_15_addr = 8'hf;
  assign ram_0_MPORT_15_mask = 1'h1;
  assign ram_0_MPORT_15_en = reset;
  assign ram_0_MPORT_16_data = 2'h0;
  assign ram_0_MPORT_16_addr = 8'h10;
  assign ram_0_MPORT_16_mask = 1'h1;
  assign ram_0_MPORT_16_en = reset;
  assign ram_0_MPORT_17_data = 2'h0;
  assign ram_0_MPORT_17_addr = 8'h11;
  assign ram_0_MPORT_17_mask = 1'h1;
  assign ram_0_MPORT_17_en = reset;
  assign ram_0_MPORT_18_data = 2'h0;
  assign ram_0_MPORT_18_addr = 8'h12;
  assign ram_0_MPORT_18_mask = 1'h1;
  assign ram_0_MPORT_18_en = reset;
  assign ram_0_MPORT_19_data = 2'h0;
  assign ram_0_MPORT_19_addr = 8'h13;
  assign ram_0_MPORT_19_mask = 1'h1;
  assign ram_0_MPORT_19_en = reset;
  assign ram_0_MPORT_20_data = 2'h0;
  assign ram_0_MPORT_20_addr = 8'h14;
  assign ram_0_MPORT_20_mask = 1'h1;
  assign ram_0_MPORT_20_en = reset;
  assign ram_0_MPORT_21_data = 2'h0;
  assign ram_0_MPORT_21_addr = 8'h15;
  assign ram_0_MPORT_21_mask = 1'h1;
  assign ram_0_MPORT_21_en = reset;
  assign ram_0_MPORT_22_data = 2'h0;
  assign ram_0_MPORT_22_addr = 8'h16;
  assign ram_0_MPORT_22_mask = 1'h1;
  assign ram_0_MPORT_22_en = reset;
  assign ram_0_MPORT_23_data = 2'h0;
  assign ram_0_MPORT_23_addr = 8'h17;
  assign ram_0_MPORT_23_mask = 1'h1;
  assign ram_0_MPORT_23_en = reset;
  assign ram_0_MPORT_24_data = 2'h0;
  assign ram_0_MPORT_24_addr = 8'h18;
  assign ram_0_MPORT_24_mask = 1'h1;
  assign ram_0_MPORT_24_en = reset;
  assign ram_0_MPORT_25_data = 2'h0;
  assign ram_0_MPORT_25_addr = 8'h19;
  assign ram_0_MPORT_25_mask = 1'h1;
  assign ram_0_MPORT_25_en = reset;
  assign ram_0_MPORT_26_data = 2'h0;
  assign ram_0_MPORT_26_addr = 8'h1a;
  assign ram_0_MPORT_26_mask = 1'h1;
  assign ram_0_MPORT_26_en = reset;
  assign ram_0_MPORT_27_data = 2'h0;
  assign ram_0_MPORT_27_addr = 8'h1b;
  assign ram_0_MPORT_27_mask = 1'h1;
  assign ram_0_MPORT_27_en = reset;
  assign ram_0_MPORT_28_data = 2'h0;
  assign ram_0_MPORT_28_addr = 8'h1c;
  assign ram_0_MPORT_28_mask = 1'h1;
  assign ram_0_MPORT_28_en = reset;
  assign ram_0_MPORT_29_data = 2'h0;
  assign ram_0_MPORT_29_addr = 8'h1d;
  assign ram_0_MPORT_29_mask = 1'h1;
  assign ram_0_MPORT_29_en = reset;
  assign ram_0_MPORT_30_data = 2'h0;
  assign ram_0_MPORT_30_addr = 8'h1e;
  assign ram_0_MPORT_30_mask = 1'h1;
  assign ram_0_MPORT_30_en = reset;
  assign ram_0_MPORT_31_data = 2'h0;
  assign ram_0_MPORT_31_addr = 8'h1f;
  assign ram_0_MPORT_31_mask = 1'h1;
  assign ram_0_MPORT_31_en = reset;
  assign ram_0_MPORT_32_data = 2'h0;
  assign ram_0_MPORT_32_addr = 8'h20;
  assign ram_0_MPORT_32_mask = 1'h1;
  assign ram_0_MPORT_32_en = reset;
  assign ram_0_MPORT_33_data = 2'h0;
  assign ram_0_MPORT_33_addr = 8'h21;
  assign ram_0_MPORT_33_mask = 1'h1;
  assign ram_0_MPORT_33_en = reset;
  assign ram_0_MPORT_34_data = 2'h0;
  assign ram_0_MPORT_34_addr = 8'h22;
  assign ram_0_MPORT_34_mask = 1'h1;
  assign ram_0_MPORT_34_en = reset;
  assign ram_0_MPORT_35_data = 2'h0;
  assign ram_0_MPORT_35_addr = 8'h23;
  assign ram_0_MPORT_35_mask = 1'h1;
  assign ram_0_MPORT_35_en = reset;
  assign ram_0_MPORT_36_data = 2'h0;
  assign ram_0_MPORT_36_addr = 8'h24;
  assign ram_0_MPORT_36_mask = 1'h1;
  assign ram_0_MPORT_36_en = reset;
  assign ram_0_MPORT_37_data = 2'h0;
  assign ram_0_MPORT_37_addr = 8'h25;
  assign ram_0_MPORT_37_mask = 1'h1;
  assign ram_0_MPORT_37_en = reset;
  assign ram_0_MPORT_38_data = 2'h0;
  assign ram_0_MPORT_38_addr = 8'h26;
  assign ram_0_MPORT_38_mask = 1'h1;
  assign ram_0_MPORT_38_en = reset;
  assign ram_0_MPORT_39_data = 2'h0;
  assign ram_0_MPORT_39_addr = 8'h27;
  assign ram_0_MPORT_39_mask = 1'h1;
  assign ram_0_MPORT_39_en = reset;
  assign ram_0_MPORT_40_data = 2'h0;
  assign ram_0_MPORT_40_addr = 8'h28;
  assign ram_0_MPORT_40_mask = 1'h1;
  assign ram_0_MPORT_40_en = reset;
  assign ram_0_MPORT_41_data = 2'h0;
  assign ram_0_MPORT_41_addr = 8'h29;
  assign ram_0_MPORT_41_mask = 1'h1;
  assign ram_0_MPORT_41_en = reset;
  assign ram_0_MPORT_42_data = 2'h0;
  assign ram_0_MPORT_42_addr = 8'h2a;
  assign ram_0_MPORT_42_mask = 1'h1;
  assign ram_0_MPORT_42_en = reset;
  assign ram_0_MPORT_43_data = 2'h0;
  assign ram_0_MPORT_43_addr = 8'h2b;
  assign ram_0_MPORT_43_mask = 1'h1;
  assign ram_0_MPORT_43_en = reset;
  assign ram_0_MPORT_44_data = 2'h0;
  assign ram_0_MPORT_44_addr = 8'h2c;
  assign ram_0_MPORT_44_mask = 1'h1;
  assign ram_0_MPORT_44_en = reset;
  assign ram_0_MPORT_45_data = 2'h0;
  assign ram_0_MPORT_45_addr = 8'h2d;
  assign ram_0_MPORT_45_mask = 1'h1;
  assign ram_0_MPORT_45_en = reset;
  assign ram_0_MPORT_46_data = 2'h0;
  assign ram_0_MPORT_46_addr = 8'h2e;
  assign ram_0_MPORT_46_mask = 1'h1;
  assign ram_0_MPORT_46_en = reset;
  assign ram_0_MPORT_47_data = 2'h0;
  assign ram_0_MPORT_47_addr = 8'h2f;
  assign ram_0_MPORT_47_mask = 1'h1;
  assign ram_0_MPORT_47_en = reset;
  assign ram_0_MPORT_48_data = 2'h0;
  assign ram_0_MPORT_48_addr = 8'h30;
  assign ram_0_MPORT_48_mask = 1'h1;
  assign ram_0_MPORT_48_en = reset;
  assign ram_0_MPORT_49_data = 2'h0;
  assign ram_0_MPORT_49_addr = 8'h31;
  assign ram_0_MPORT_49_mask = 1'h1;
  assign ram_0_MPORT_49_en = reset;
  assign ram_0_MPORT_50_data = 2'h0;
  assign ram_0_MPORT_50_addr = 8'h32;
  assign ram_0_MPORT_50_mask = 1'h1;
  assign ram_0_MPORT_50_en = reset;
  assign ram_0_MPORT_51_data = 2'h0;
  assign ram_0_MPORT_51_addr = 8'h33;
  assign ram_0_MPORT_51_mask = 1'h1;
  assign ram_0_MPORT_51_en = reset;
  assign ram_0_MPORT_52_data = 2'h0;
  assign ram_0_MPORT_52_addr = 8'h34;
  assign ram_0_MPORT_52_mask = 1'h1;
  assign ram_0_MPORT_52_en = reset;
  assign ram_0_MPORT_53_data = 2'h0;
  assign ram_0_MPORT_53_addr = 8'h35;
  assign ram_0_MPORT_53_mask = 1'h1;
  assign ram_0_MPORT_53_en = reset;
  assign ram_0_MPORT_54_data = 2'h0;
  assign ram_0_MPORT_54_addr = 8'h36;
  assign ram_0_MPORT_54_mask = 1'h1;
  assign ram_0_MPORT_54_en = reset;
  assign ram_0_MPORT_55_data = 2'h0;
  assign ram_0_MPORT_55_addr = 8'h37;
  assign ram_0_MPORT_55_mask = 1'h1;
  assign ram_0_MPORT_55_en = reset;
  assign ram_0_MPORT_56_data = 2'h0;
  assign ram_0_MPORT_56_addr = 8'h38;
  assign ram_0_MPORT_56_mask = 1'h1;
  assign ram_0_MPORT_56_en = reset;
  assign ram_0_MPORT_57_data = 2'h0;
  assign ram_0_MPORT_57_addr = 8'h39;
  assign ram_0_MPORT_57_mask = 1'h1;
  assign ram_0_MPORT_57_en = reset;
  assign ram_0_MPORT_58_data = 2'h0;
  assign ram_0_MPORT_58_addr = 8'h3a;
  assign ram_0_MPORT_58_mask = 1'h1;
  assign ram_0_MPORT_58_en = reset;
  assign ram_0_MPORT_59_data = 2'h0;
  assign ram_0_MPORT_59_addr = 8'h3b;
  assign ram_0_MPORT_59_mask = 1'h1;
  assign ram_0_MPORT_59_en = reset;
  assign ram_0_MPORT_60_data = 2'h0;
  assign ram_0_MPORT_60_addr = 8'h3c;
  assign ram_0_MPORT_60_mask = 1'h1;
  assign ram_0_MPORT_60_en = reset;
  assign ram_0_MPORT_61_data = 2'h0;
  assign ram_0_MPORT_61_addr = 8'h3d;
  assign ram_0_MPORT_61_mask = 1'h1;
  assign ram_0_MPORT_61_en = reset;
  assign ram_0_MPORT_62_data = 2'h0;
  assign ram_0_MPORT_62_addr = 8'h3e;
  assign ram_0_MPORT_62_mask = 1'h1;
  assign ram_0_MPORT_62_en = reset;
  assign ram_0_MPORT_63_data = 2'h0;
  assign ram_0_MPORT_63_addr = 8'h3f;
  assign ram_0_MPORT_63_mask = 1'h1;
  assign ram_0_MPORT_63_en = reset;
  assign ram_0_MPORT_64_data = 2'h0;
  assign ram_0_MPORT_64_addr = 8'h40;
  assign ram_0_MPORT_64_mask = 1'h1;
  assign ram_0_MPORT_64_en = reset;
  assign ram_0_MPORT_65_data = 2'h0;
  assign ram_0_MPORT_65_addr = 8'h41;
  assign ram_0_MPORT_65_mask = 1'h1;
  assign ram_0_MPORT_65_en = reset;
  assign ram_0_MPORT_66_data = 2'h0;
  assign ram_0_MPORT_66_addr = 8'h42;
  assign ram_0_MPORT_66_mask = 1'h1;
  assign ram_0_MPORT_66_en = reset;
  assign ram_0_MPORT_67_data = 2'h0;
  assign ram_0_MPORT_67_addr = 8'h43;
  assign ram_0_MPORT_67_mask = 1'h1;
  assign ram_0_MPORT_67_en = reset;
  assign ram_0_MPORT_68_data = 2'h0;
  assign ram_0_MPORT_68_addr = 8'h44;
  assign ram_0_MPORT_68_mask = 1'h1;
  assign ram_0_MPORT_68_en = reset;
  assign ram_0_MPORT_69_data = 2'h0;
  assign ram_0_MPORT_69_addr = 8'h45;
  assign ram_0_MPORT_69_mask = 1'h1;
  assign ram_0_MPORT_69_en = reset;
  assign ram_0_MPORT_70_data = 2'h0;
  assign ram_0_MPORT_70_addr = 8'h46;
  assign ram_0_MPORT_70_mask = 1'h1;
  assign ram_0_MPORT_70_en = reset;
  assign ram_0_MPORT_71_data = 2'h0;
  assign ram_0_MPORT_71_addr = 8'h47;
  assign ram_0_MPORT_71_mask = 1'h1;
  assign ram_0_MPORT_71_en = reset;
  assign ram_0_MPORT_72_data = 2'h0;
  assign ram_0_MPORT_72_addr = 8'h48;
  assign ram_0_MPORT_72_mask = 1'h1;
  assign ram_0_MPORT_72_en = reset;
  assign ram_0_MPORT_73_data = 2'h0;
  assign ram_0_MPORT_73_addr = 8'h49;
  assign ram_0_MPORT_73_mask = 1'h1;
  assign ram_0_MPORT_73_en = reset;
  assign ram_0_MPORT_74_data = 2'h0;
  assign ram_0_MPORT_74_addr = 8'h4a;
  assign ram_0_MPORT_74_mask = 1'h1;
  assign ram_0_MPORT_74_en = reset;
  assign ram_0_MPORT_75_data = 2'h0;
  assign ram_0_MPORT_75_addr = 8'h4b;
  assign ram_0_MPORT_75_mask = 1'h1;
  assign ram_0_MPORT_75_en = reset;
  assign ram_0_MPORT_76_data = 2'h0;
  assign ram_0_MPORT_76_addr = 8'h4c;
  assign ram_0_MPORT_76_mask = 1'h1;
  assign ram_0_MPORT_76_en = reset;
  assign ram_0_MPORT_77_data = 2'h0;
  assign ram_0_MPORT_77_addr = 8'h4d;
  assign ram_0_MPORT_77_mask = 1'h1;
  assign ram_0_MPORT_77_en = reset;
  assign ram_0_MPORT_78_data = 2'h0;
  assign ram_0_MPORT_78_addr = 8'h4e;
  assign ram_0_MPORT_78_mask = 1'h1;
  assign ram_0_MPORT_78_en = reset;
  assign ram_0_MPORT_79_data = 2'h0;
  assign ram_0_MPORT_79_addr = 8'h4f;
  assign ram_0_MPORT_79_mask = 1'h1;
  assign ram_0_MPORT_79_en = reset;
  assign ram_0_MPORT_80_data = 2'h0;
  assign ram_0_MPORT_80_addr = 8'h50;
  assign ram_0_MPORT_80_mask = 1'h1;
  assign ram_0_MPORT_80_en = reset;
  assign ram_0_MPORT_81_data = 2'h0;
  assign ram_0_MPORT_81_addr = 8'h51;
  assign ram_0_MPORT_81_mask = 1'h1;
  assign ram_0_MPORT_81_en = reset;
  assign ram_0_MPORT_82_data = 2'h0;
  assign ram_0_MPORT_82_addr = 8'h52;
  assign ram_0_MPORT_82_mask = 1'h1;
  assign ram_0_MPORT_82_en = reset;
  assign ram_0_MPORT_83_data = 2'h0;
  assign ram_0_MPORT_83_addr = 8'h53;
  assign ram_0_MPORT_83_mask = 1'h1;
  assign ram_0_MPORT_83_en = reset;
  assign ram_0_MPORT_84_data = 2'h0;
  assign ram_0_MPORT_84_addr = 8'h54;
  assign ram_0_MPORT_84_mask = 1'h1;
  assign ram_0_MPORT_84_en = reset;
  assign ram_0_MPORT_85_data = 2'h0;
  assign ram_0_MPORT_85_addr = 8'h55;
  assign ram_0_MPORT_85_mask = 1'h1;
  assign ram_0_MPORT_85_en = reset;
  assign ram_0_MPORT_86_data = 2'h0;
  assign ram_0_MPORT_86_addr = 8'h56;
  assign ram_0_MPORT_86_mask = 1'h1;
  assign ram_0_MPORT_86_en = reset;
  assign ram_0_MPORT_87_data = 2'h0;
  assign ram_0_MPORT_87_addr = 8'h57;
  assign ram_0_MPORT_87_mask = 1'h1;
  assign ram_0_MPORT_87_en = reset;
  assign ram_0_MPORT_88_data = 2'h0;
  assign ram_0_MPORT_88_addr = 8'h58;
  assign ram_0_MPORT_88_mask = 1'h1;
  assign ram_0_MPORT_88_en = reset;
  assign ram_0_MPORT_89_data = 2'h0;
  assign ram_0_MPORT_89_addr = 8'h59;
  assign ram_0_MPORT_89_mask = 1'h1;
  assign ram_0_MPORT_89_en = reset;
  assign ram_0_MPORT_90_data = 2'h0;
  assign ram_0_MPORT_90_addr = 8'h5a;
  assign ram_0_MPORT_90_mask = 1'h1;
  assign ram_0_MPORT_90_en = reset;
  assign ram_0_MPORT_91_data = 2'h0;
  assign ram_0_MPORT_91_addr = 8'h5b;
  assign ram_0_MPORT_91_mask = 1'h1;
  assign ram_0_MPORT_91_en = reset;
  assign ram_0_MPORT_92_data = 2'h0;
  assign ram_0_MPORT_92_addr = 8'h5c;
  assign ram_0_MPORT_92_mask = 1'h1;
  assign ram_0_MPORT_92_en = reset;
  assign ram_0_MPORT_93_data = 2'h0;
  assign ram_0_MPORT_93_addr = 8'h5d;
  assign ram_0_MPORT_93_mask = 1'h1;
  assign ram_0_MPORT_93_en = reset;
  assign ram_0_MPORT_94_data = 2'h0;
  assign ram_0_MPORT_94_addr = 8'h5e;
  assign ram_0_MPORT_94_mask = 1'h1;
  assign ram_0_MPORT_94_en = reset;
  assign ram_0_MPORT_95_data = 2'h0;
  assign ram_0_MPORT_95_addr = 8'h5f;
  assign ram_0_MPORT_95_mask = 1'h1;
  assign ram_0_MPORT_95_en = reset;
  assign ram_0_MPORT_96_data = 2'h0;
  assign ram_0_MPORT_96_addr = 8'h60;
  assign ram_0_MPORT_96_mask = 1'h1;
  assign ram_0_MPORT_96_en = reset;
  assign ram_0_MPORT_97_data = 2'h0;
  assign ram_0_MPORT_97_addr = 8'h61;
  assign ram_0_MPORT_97_mask = 1'h1;
  assign ram_0_MPORT_97_en = reset;
  assign ram_0_MPORT_98_data = 2'h0;
  assign ram_0_MPORT_98_addr = 8'h62;
  assign ram_0_MPORT_98_mask = 1'h1;
  assign ram_0_MPORT_98_en = reset;
  assign ram_0_MPORT_99_data = 2'h0;
  assign ram_0_MPORT_99_addr = 8'h63;
  assign ram_0_MPORT_99_mask = 1'h1;
  assign ram_0_MPORT_99_en = reset;
  assign ram_0_MPORT_100_data = 2'h0;
  assign ram_0_MPORT_100_addr = 8'h64;
  assign ram_0_MPORT_100_mask = 1'h1;
  assign ram_0_MPORT_100_en = reset;
  assign ram_0_MPORT_101_data = 2'h0;
  assign ram_0_MPORT_101_addr = 8'h65;
  assign ram_0_MPORT_101_mask = 1'h1;
  assign ram_0_MPORT_101_en = reset;
  assign ram_0_MPORT_102_data = 2'h0;
  assign ram_0_MPORT_102_addr = 8'h66;
  assign ram_0_MPORT_102_mask = 1'h1;
  assign ram_0_MPORT_102_en = reset;
  assign ram_0_MPORT_103_data = 2'h0;
  assign ram_0_MPORT_103_addr = 8'h67;
  assign ram_0_MPORT_103_mask = 1'h1;
  assign ram_0_MPORT_103_en = reset;
  assign ram_0_MPORT_104_data = 2'h0;
  assign ram_0_MPORT_104_addr = 8'h68;
  assign ram_0_MPORT_104_mask = 1'h1;
  assign ram_0_MPORT_104_en = reset;
  assign ram_0_MPORT_105_data = 2'h0;
  assign ram_0_MPORT_105_addr = 8'h69;
  assign ram_0_MPORT_105_mask = 1'h1;
  assign ram_0_MPORT_105_en = reset;
  assign ram_0_MPORT_106_data = 2'h0;
  assign ram_0_MPORT_106_addr = 8'h6a;
  assign ram_0_MPORT_106_mask = 1'h1;
  assign ram_0_MPORT_106_en = reset;
  assign ram_0_MPORT_107_data = 2'h0;
  assign ram_0_MPORT_107_addr = 8'h6b;
  assign ram_0_MPORT_107_mask = 1'h1;
  assign ram_0_MPORT_107_en = reset;
  assign ram_0_MPORT_108_data = 2'h0;
  assign ram_0_MPORT_108_addr = 8'h6c;
  assign ram_0_MPORT_108_mask = 1'h1;
  assign ram_0_MPORT_108_en = reset;
  assign ram_0_MPORT_109_data = 2'h0;
  assign ram_0_MPORT_109_addr = 8'h6d;
  assign ram_0_MPORT_109_mask = 1'h1;
  assign ram_0_MPORT_109_en = reset;
  assign ram_0_MPORT_110_data = 2'h0;
  assign ram_0_MPORT_110_addr = 8'h6e;
  assign ram_0_MPORT_110_mask = 1'h1;
  assign ram_0_MPORT_110_en = reset;
  assign ram_0_MPORT_111_data = 2'h0;
  assign ram_0_MPORT_111_addr = 8'h6f;
  assign ram_0_MPORT_111_mask = 1'h1;
  assign ram_0_MPORT_111_en = reset;
  assign ram_0_MPORT_112_data = 2'h0;
  assign ram_0_MPORT_112_addr = 8'h70;
  assign ram_0_MPORT_112_mask = 1'h1;
  assign ram_0_MPORT_112_en = reset;
  assign ram_0_MPORT_113_data = 2'h0;
  assign ram_0_MPORT_113_addr = 8'h71;
  assign ram_0_MPORT_113_mask = 1'h1;
  assign ram_0_MPORT_113_en = reset;
  assign ram_0_MPORT_114_data = 2'h0;
  assign ram_0_MPORT_114_addr = 8'h72;
  assign ram_0_MPORT_114_mask = 1'h1;
  assign ram_0_MPORT_114_en = reset;
  assign ram_0_MPORT_115_data = 2'h0;
  assign ram_0_MPORT_115_addr = 8'h73;
  assign ram_0_MPORT_115_mask = 1'h1;
  assign ram_0_MPORT_115_en = reset;
  assign ram_0_MPORT_116_data = 2'h0;
  assign ram_0_MPORT_116_addr = 8'h74;
  assign ram_0_MPORT_116_mask = 1'h1;
  assign ram_0_MPORT_116_en = reset;
  assign ram_0_MPORT_117_data = 2'h0;
  assign ram_0_MPORT_117_addr = 8'h75;
  assign ram_0_MPORT_117_mask = 1'h1;
  assign ram_0_MPORT_117_en = reset;
  assign ram_0_MPORT_118_data = 2'h0;
  assign ram_0_MPORT_118_addr = 8'h76;
  assign ram_0_MPORT_118_mask = 1'h1;
  assign ram_0_MPORT_118_en = reset;
  assign ram_0_MPORT_119_data = 2'h0;
  assign ram_0_MPORT_119_addr = 8'h77;
  assign ram_0_MPORT_119_mask = 1'h1;
  assign ram_0_MPORT_119_en = reset;
  assign ram_0_MPORT_120_data = 2'h0;
  assign ram_0_MPORT_120_addr = 8'h78;
  assign ram_0_MPORT_120_mask = 1'h1;
  assign ram_0_MPORT_120_en = reset;
  assign ram_0_MPORT_121_data = 2'h0;
  assign ram_0_MPORT_121_addr = 8'h79;
  assign ram_0_MPORT_121_mask = 1'h1;
  assign ram_0_MPORT_121_en = reset;
  assign ram_0_MPORT_122_data = 2'h0;
  assign ram_0_MPORT_122_addr = 8'h7a;
  assign ram_0_MPORT_122_mask = 1'h1;
  assign ram_0_MPORT_122_en = reset;
  assign ram_0_MPORT_123_data = 2'h0;
  assign ram_0_MPORT_123_addr = 8'h7b;
  assign ram_0_MPORT_123_mask = 1'h1;
  assign ram_0_MPORT_123_en = reset;
  assign ram_0_MPORT_124_data = 2'h0;
  assign ram_0_MPORT_124_addr = 8'h7c;
  assign ram_0_MPORT_124_mask = 1'h1;
  assign ram_0_MPORT_124_en = reset;
  assign ram_0_MPORT_125_data = 2'h0;
  assign ram_0_MPORT_125_addr = 8'h7d;
  assign ram_0_MPORT_125_mask = 1'h1;
  assign ram_0_MPORT_125_en = reset;
  assign ram_0_MPORT_126_data = 2'h0;
  assign ram_0_MPORT_126_addr = 8'h7e;
  assign ram_0_MPORT_126_mask = 1'h1;
  assign ram_0_MPORT_126_en = reset;
  assign ram_0_MPORT_127_data = 2'h0;
  assign ram_0_MPORT_127_addr = 8'h7f;
  assign ram_0_MPORT_127_mask = 1'h1;
  assign ram_0_MPORT_127_en = reset;
  assign ram_0_MPORT_128_data = 2'h0;
  assign ram_0_MPORT_128_addr = 8'h80;
  assign ram_0_MPORT_128_mask = 1'h1;
  assign ram_0_MPORT_128_en = reset;
  assign ram_0_MPORT_129_data = 2'h0;
  assign ram_0_MPORT_129_addr = 8'h81;
  assign ram_0_MPORT_129_mask = 1'h1;
  assign ram_0_MPORT_129_en = reset;
  assign ram_0_MPORT_130_data = 2'h0;
  assign ram_0_MPORT_130_addr = 8'h82;
  assign ram_0_MPORT_130_mask = 1'h1;
  assign ram_0_MPORT_130_en = reset;
  assign ram_0_MPORT_131_data = 2'h0;
  assign ram_0_MPORT_131_addr = 8'h83;
  assign ram_0_MPORT_131_mask = 1'h1;
  assign ram_0_MPORT_131_en = reset;
  assign ram_0_MPORT_132_data = 2'h0;
  assign ram_0_MPORT_132_addr = 8'h84;
  assign ram_0_MPORT_132_mask = 1'h1;
  assign ram_0_MPORT_132_en = reset;
  assign ram_0_MPORT_133_data = 2'h0;
  assign ram_0_MPORT_133_addr = 8'h85;
  assign ram_0_MPORT_133_mask = 1'h1;
  assign ram_0_MPORT_133_en = reset;
  assign ram_0_MPORT_134_data = 2'h0;
  assign ram_0_MPORT_134_addr = 8'h86;
  assign ram_0_MPORT_134_mask = 1'h1;
  assign ram_0_MPORT_134_en = reset;
  assign ram_0_MPORT_135_data = 2'h0;
  assign ram_0_MPORT_135_addr = 8'h87;
  assign ram_0_MPORT_135_mask = 1'h1;
  assign ram_0_MPORT_135_en = reset;
  assign ram_0_MPORT_136_data = 2'h0;
  assign ram_0_MPORT_136_addr = 8'h88;
  assign ram_0_MPORT_136_mask = 1'h1;
  assign ram_0_MPORT_136_en = reset;
  assign ram_0_MPORT_137_data = 2'h0;
  assign ram_0_MPORT_137_addr = 8'h89;
  assign ram_0_MPORT_137_mask = 1'h1;
  assign ram_0_MPORT_137_en = reset;
  assign ram_0_MPORT_138_data = 2'h0;
  assign ram_0_MPORT_138_addr = 8'h8a;
  assign ram_0_MPORT_138_mask = 1'h1;
  assign ram_0_MPORT_138_en = reset;
  assign ram_0_MPORT_139_data = 2'h0;
  assign ram_0_MPORT_139_addr = 8'h8b;
  assign ram_0_MPORT_139_mask = 1'h1;
  assign ram_0_MPORT_139_en = reset;
  assign ram_0_MPORT_140_data = 2'h0;
  assign ram_0_MPORT_140_addr = 8'h8c;
  assign ram_0_MPORT_140_mask = 1'h1;
  assign ram_0_MPORT_140_en = reset;
  assign ram_0_MPORT_141_data = 2'h0;
  assign ram_0_MPORT_141_addr = 8'h8d;
  assign ram_0_MPORT_141_mask = 1'h1;
  assign ram_0_MPORT_141_en = reset;
  assign ram_0_MPORT_142_data = 2'h0;
  assign ram_0_MPORT_142_addr = 8'h8e;
  assign ram_0_MPORT_142_mask = 1'h1;
  assign ram_0_MPORT_142_en = reset;
  assign ram_0_MPORT_143_data = 2'h0;
  assign ram_0_MPORT_143_addr = 8'h8f;
  assign ram_0_MPORT_143_mask = 1'h1;
  assign ram_0_MPORT_143_en = reset;
  assign ram_0_MPORT_144_data = 2'h0;
  assign ram_0_MPORT_144_addr = 8'h90;
  assign ram_0_MPORT_144_mask = 1'h1;
  assign ram_0_MPORT_144_en = reset;
  assign ram_0_MPORT_145_data = 2'h0;
  assign ram_0_MPORT_145_addr = 8'h91;
  assign ram_0_MPORT_145_mask = 1'h1;
  assign ram_0_MPORT_145_en = reset;
  assign ram_0_MPORT_146_data = 2'h0;
  assign ram_0_MPORT_146_addr = 8'h92;
  assign ram_0_MPORT_146_mask = 1'h1;
  assign ram_0_MPORT_146_en = reset;
  assign ram_0_MPORT_147_data = 2'h0;
  assign ram_0_MPORT_147_addr = 8'h93;
  assign ram_0_MPORT_147_mask = 1'h1;
  assign ram_0_MPORT_147_en = reset;
  assign ram_0_MPORT_148_data = 2'h0;
  assign ram_0_MPORT_148_addr = 8'h94;
  assign ram_0_MPORT_148_mask = 1'h1;
  assign ram_0_MPORT_148_en = reset;
  assign ram_0_MPORT_149_data = 2'h0;
  assign ram_0_MPORT_149_addr = 8'h95;
  assign ram_0_MPORT_149_mask = 1'h1;
  assign ram_0_MPORT_149_en = reset;
  assign ram_0_MPORT_150_data = 2'h0;
  assign ram_0_MPORT_150_addr = 8'h96;
  assign ram_0_MPORT_150_mask = 1'h1;
  assign ram_0_MPORT_150_en = reset;
  assign ram_0_MPORT_151_data = 2'h0;
  assign ram_0_MPORT_151_addr = 8'h97;
  assign ram_0_MPORT_151_mask = 1'h1;
  assign ram_0_MPORT_151_en = reset;
  assign ram_0_MPORT_152_data = 2'h0;
  assign ram_0_MPORT_152_addr = 8'h98;
  assign ram_0_MPORT_152_mask = 1'h1;
  assign ram_0_MPORT_152_en = reset;
  assign ram_0_MPORT_153_data = 2'h0;
  assign ram_0_MPORT_153_addr = 8'h99;
  assign ram_0_MPORT_153_mask = 1'h1;
  assign ram_0_MPORT_153_en = reset;
  assign ram_0_MPORT_154_data = 2'h0;
  assign ram_0_MPORT_154_addr = 8'h9a;
  assign ram_0_MPORT_154_mask = 1'h1;
  assign ram_0_MPORT_154_en = reset;
  assign ram_0_MPORT_155_data = 2'h0;
  assign ram_0_MPORT_155_addr = 8'h9b;
  assign ram_0_MPORT_155_mask = 1'h1;
  assign ram_0_MPORT_155_en = reset;
  assign ram_0_MPORT_156_data = 2'h0;
  assign ram_0_MPORT_156_addr = 8'h9c;
  assign ram_0_MPORT_156_mask = 1'h1;
  assign ram_0_MPORT_156_en = reset;
  assign ram_0_MPORT_157_data = 2'h0;
  assign ram_0_MPORT_157_addr = 8'h9d;
  assign ram_0_MPORT_157_mask = 1'h1;
  assign ram_0_MPORT_157_en = reset;
  assign ram_0_MPORT_158_data = 2'h0;
  assign ram_0_MPORT_158_addr = 8'h9e;
  assign ram_0_MPORT_158_mask = 1'h1;
  assign ram_0_MPORT_158_en = reset;
  assign ram_0_MPORT_159_data = 2'h0;
  assign ram_0_MPORT_159_addr = 8'h9f;
  assign ram_0_MPORT_159_mask = 1'h1;
  assign ram_0_MPORT_159_en = reset;
  assign ram_0_MPORT_160_data = 2'h0;
  assign ram_0_MPORT_160_addr = 8'ha0;
  assign ram_0_MPORT_160_mask = 1'h1;
  assign ram_0_MPORT_160_en = reset;
  assign ram_0_MPORT_161_data = 2'h0;
  assign ram_0_MPORT_161_addr = 8'ha1;
  assign ram_0_MPORT_161_mask = 1'h1;
  assign ram_0_MPORT_161_en = reset;
  assign ram_0_MPORT_162_data = 2'h0;
  assign ram_0_MPORT_162_addr = 8'ha2;
  assign ram_0_MPORT_162_mask = 1'h1;
  assign ram_0_MPORT_162_en = reset;
  assign ram_0_MPORT_163_data = 2'h0;
  assign ram_0_MPORT_163_addr = 8'ha3;
  assign ram_0_MPORT_163_mask = 1'h1;
  assign ram_0_MPORT_163_en = reset;
  assign ram_0_MPORT_164_data = 2'h0;
  assign ram_0_MPORT_164_addr = 8'ha4;
  assign ram_0_MPORT_164_mask = 1'h1;
  assign ram_0_MPORT_164_en = reset;
  assign ram_0_MPORT_165_data = 2'h0;
  assign ram_0_MPORT_165_addr = 8'ha5;
  assign ram_0_MPORT_165_mask = 1'h1;
  assign ram_0_MPORT_165_en = reset;
  assign ram_0_MPORT_166_data = 2'h0;
  assign ram_0_MPORT_166_addr = 8'ha6;
  assign ram_0_MPORT_166_mask = 1'h1;
  assign ram_0_MPORT_166_en = reset;
  assign ram_0_MPORT_167_data = 2'h0;
  assign ram_0_MPORT_167_addr = 8'ha7;
  assign ram_0_MPORT_167_mask = 1'h1;
  assign ram_0_MPORT_167_en = reset;
  assign ram_0_MPORT_168_data = 2'h0;
  assign ram_0_MPORT_168_addr = 8'ha8;
  assign ram_0_MPORT_168_mask = 1'h1;
  assign ram_0_MPORT_168_en = reset;
  assign ram_0_MPORT_169_data = 2'h0;
  assign ram_0_MPORT_169_addr = 8'ha9;
  assign ram_0_MPORT_169_mask = 1'h1;
  assign ram_0_MPORT_169_en = reset;
  assign ram_0_MPORT_170_data = 2'h0;
  assign ram_0_MPORT_170_addr = 8'haa;
  assign ram_0_MPORT_170_mask = 1'h1;
  assign ram_0_MPORT_170_en = reset;
  assign ram_0_MPORT_171_data = 2'h0;
  assign ram_0_MPORT_171_addr = 8'hab;
  assign ram_0_MPORT_171_mask = 1'h1;
  assign ram_0_MPORT_171_en = reset;
  assign ram_0_MPORT_172_data = 2'h0;
  assign ram_0_MPORT_172_addr = 8'hac;
  assign ram_0_MPORT_172_mask = 1'h1;
  assign ram_0_MPORT_172_en = reset;
  assign ram_0_MPORT_173_data = 2'h0;
  assign ram_0_MPORT_173_addr = 8'had;
  assign ram_0_MPORT_173_mask = 1'h1;
  assign ram_0_MPORT_173_en = reset;
  assign ram_0_MPORT_174_data = 2'h0;
  assign ram_0_MPORT_174_addr = 8'hae;
  assign ram_0_MPORT_174_mask = 1'h1;
  assign ram_0_MPORT_174_en = reset;
  assign ram_0_MPORT_175_data = 2'h0;
  assign ram_0_MPORT_175_addr = 8'haf;
  assign ram_0_MPORT_175_mask = 1'h1;
  assign ram_0_MPORT_175_en = reset;
  assign ram_0_MPORT_176_data = 2'h0;
  assign ram_0_MPORT_176_addr = 8'hb0;
  assign ram_0_MPORT_176_mask = 1'h1;
  assign ram_0_MPORT_176_en = reset;
  assign ram_0_MPORT_177_data = 2'h0;
  assign ram_0_MPORT_177_addr = 8'hb1;
  assign ram_0_MPORT_177_mask = 1'h1;
  assign ram_0_MPORT_177_en = reset;
  assign ram_0_MPORT_178_data = 2'h0;
  assign ram_0_MPORT_178_addr = 8'hb2;
  assign ram_0_MPORT_178_mask = 1'h1;
  assign ram_0_MPORT_178_en = reset;
  assign ram_0_MPORT_179_data = 2'h0;
  assign ram_0_MPORT_179_addr = 8'hb3;
  assign ram_0_MPORT_179_mask = 1'h1;
  assign ram_0_MPORT_179_en = reset;
  assign ram_0_MPORT_180_data = 2'h0;
  assign ram_0_MPORT_180_addr = 8'hb4;
  assign ram_0_MPORT_180_mask = 1'h1;
  assign ram_0_MPORT_180_en = reset;
  assign ram_0_MPORT_181_data = 2'h0;
  assign ram_0_MPORT_181_addr = 8'hb5;
  assign ram_0_MPORT_181_mask = 1'h1;
  assign ram_0_MPORT_181_en = reset;
  assign ram_0_MPORT_182_data = 2'h0;
  assign ram_0_MPORT_182_addr = 8'hb6;
  assign ram_0_MPORT_182_mask = 1'h1;
  assign ram_0_MPORT_182_en = reset;
  assign ram_0_MPORT_183_data = 2'h0;
  assign ram_0_MPORT_183_addr = 8'hb7;
  assign ram_0_MPORT_183_mask = 1'h1;
  assign ram_0_MPORT_183_en = reset;
  assign ram_0_MPORT_184_data = 2'h0;
  assign ram_0_MPORT_184_addr = 8'hb8;
  assign ram_0_MPORT_184_mask = 1'h1;
  assign ram_0_MPORT_184_en = reset;
  assign ram_0_MPORT_185_data = 2'h0;
  assign ram_0_MPORT_185_addr = 8'hb9;
  assign ram_0_MPORT_185_mask = 1'h1;
  assign ram_0_MPORT_185_en = reset;
  assign ram_0_MPORT_186_data = 2'h0;
  assign ram_0_MPORT_186_addr = 8'hba;
  assign ram_0_MPORT_186_mask = 1'h1;
  assign ram_0_MPORT_186_en = reset;
  assign ram_0_MPORT_187_data = 2'h0;
  assign ram_0_MPORT_187_addr = 8'hbb;
  assign ram_0_MPORT_187_mask = 1'h1;
  assign ram_0_MPORT_187_en = reset;
  assign ram_0_MPORT_188_data = 2'h0;
  assign ram_0_MPORT_188_addr = 8'hbc;
  assign ram_0_MPORT_188_mask = 1'h1;
  assign ram_0_MPORT_188_en = reset;
  assign ram_0_MPORT_189_data = 2'h0;
  assign ram_0_MPORT_189_addr = 8'hbd;
  assign ram_0_MPORT_189_mask = 1'h1;
  assign ram_0_MPORT_189_en = reset;
  assign ram_0_MPORT_190_data = 2'h0;
  assign ram_0_MPORT_190_addr = 8'hbe;
  assign ram_0_MPORT_190_mask = 1'h1;
  assign ram_0_MPORT_190_en = reset;
  assign ram_0_MPORT_191_data = 2'h0;
  assign ram_0_MPORT_191_addr = 8'hbf;
  assign ram_0_MPORT_191_mask = 1'h1;
  assign ram_0_MPORT_191_en = reset;
  assign ram_0_MPORT_192_data = 2'h0;
  assign ram_0_MPORT_192_addr = 8'hc0;
  assign ram_0_MPORT_192_mask = 1'h1;
  assign ram_0_MPORT_192_en = reset;
  assign ram_0_MPORT_193_data = 2'h0;
  assign ram_0_MPORT_193_addr = 8'hc1;
  assign ram_0_MPORT_193_mask = 1'h1;
  assign ram_0_MPORT_193_en = reset;
  assign ram_0_MPORT_194_data = 2'h0;
  assign ram_0_MPORT_194_addr = 8'hc2;
  assign ram_0_MPORT_194_mask = 1'h1;
  assign ram_0_MPORT_194_en = reset;
  assign ram_0_MPORT_195_data = 2'h0;
  assign ram_0_MPORT_195_addr = 8'hc3;
  assign ram_0_MPORT_195_mask = 1'h1;
  assign ram_0_MPORT_195_en = reset;
  assign ram_0_MPORT_196_data = 2'h0;
  assign ram_0_MPORT_196_addr = 8'hc4;
  assign ram_0_MPORT_196_mask = 1'h1;
  assign ram_0_MPORT_196_en = reset;
  assign ram_0_MPORT_197_data = 2'h0;
  assign ram_0_MPORT_197_addr = 8'hc5;
  assign ram_0_MPORT_197_mask = 1'h1;
  assign ram_0_MPORT_197_en = reset;
  assign ram_0_MPORT_198_data = 2'h0;
  assign ram_0_MPORT_198_addr = 8'hc6;
  assign ram_0_MPORT_198_mask = 1'h1;
  assign ram_0_MPORT_198_en = reset;
  assign ram_0_MPORT_199_data = 2'h0;
  assign ram_0_MPORT_199_addr = 8'hc7;
  assign ram_0_MPORT_199_mask = 1'h1;
  assign ram_0_MPORT_199_en = reset;
  assign ram_0_MPORT_200_data = 2'h0;
  assign ram_0_MPORT_200_addr = 8'hc8;
  assign ram_0_MPORT_200_mask = 1'h1;
  assign ram_0_MPORT_200_en = reset;
  assign ram_0_MPORT_201_data = 2'h0;
  assign ram_0_MPORT_201_addr = 8'hc9;
  assign ram_0_MPORT_201_mask = 1'h1;
  assign ram_0_MPORT_201_en = reset;
  assign ram_0_MPORT_202_data = 2'h0;
  assign ram_0_MPORT_202_addr = 8'hca;
  assign ram_0_MPORT_202_mask = 1'h1;
  assign ram_0_MPORT_202_en = reset;
  assign ram_0_MPORT_203_data = 2'h0;
  assign ram_0_MPORT_203_addr = 8'hcb;
  assign ram_0_MPORT_203_mask = 1'h1;
  assign ram_0_MPORT_203_en = reset;
  assign ram_0_MPORT_204_data = 2'h0;
  assign ram_0_MPORT_204_addr = 8'hcc;
  assign ram_0_MPORT_204_mask = 1'h1;
  assign ram_0_MPORT_204_en = reset;
  assign ram_0_MPORT_205_data = 2'h0;
  assign ram_0_MPORT_205_addr = 8'hcd;
  assign ram_0_MPORT_205_mask = 1'h1;
  assign ram_0_MPORT_205_en = reset;
  assign ram_0_MPORT_206_data = 2'h0;
  assign ram_0_MPORT_206_addr = 8'hce;
  assign ram_0_MPORT_206_mask = 1'h1;
  assign ram_0_MPORT_206_en = reset;
  assign ram_0_MPORT_207_data = 2'h0;
  assign ram_0_MPORT_207_addr = 8'hcf;
  assign ram_0_MPORT_207_mask = 1'h1;
  assign ram_0_MPORT_207_en = reset;
  assign ram_0_MPORT_208_data = 2'h0;
  assign ram_0_MPORT_208_addr = 8'hd0;
  assign ram_0_MPORT_208_mask = 1'h1;
  assign ram_0_MPORT_208_en = reset;
  assign ram_0_MPORT_209_data = 2'h0;
  assign ram_0_MPORT_209_addr = 8'hd1;
  assign ram_0_MPORT_209_mask = 1'h1;
  assign ram_0_MPORT_209_en = reset;
  assign ram_0_MPORT_210_data = 2'h0;
  assign ram_0_MPORT_210_addr = 8'hd2;
  assign ram_0_MPORT_210_mask = 1'h1;
  assign ram_0_MPORT_210_en = reset;
  assign ram_0_MPORT_211_data = 2'h0;
  assign ram_0_MPORT_211_addr = 8'hd3;
  assign ram_0_MPORT_211_mask = 1'h1;
  assign ram_0_MPORT_211_en = reset;
  assign ram_0_MPORT_212_data = 2'h0;
  assign ram_0_MPORT_212_addr = 8'hd4;
  assign ram_0_MPORT_212_mask = 1'h1;
  assign ram_0_MPORT_212_en = reset;
  assign ram_0_MPORT_213_data = 2'h0;
  assign ram_0_MPORT_213_addr = 8'hd5;
  assign ram_0_MPORT_213_mask = 1'h1;
  assign ram_0_MPORT_213_en = reset;
  assign ram_0_MPORT_214_data = 2'h0;
  assign ram_0_MPORT_214_addr = 8'hd6;
  assign ram_0_MPORT_214_mask = 1'h1;
  assign ram_0_MPORT_214_en = reset;
  assign ram_0_MPORT_215_data = 2'h0;
  assign ram_0_MPORT_215_addr = 8'hd7;
  assign ram_0_MPORT_215_mask = 1'h1;
  assign ram_0_MPORT_215_en = reset;
  assign ram_0_MPORT_216_data = 2'h0;
  assign ram_0_MPORT_216_addr = 8'hd8;
  assign ram_0_MPORT_216_mask = 1'h1;
  assign ram_0_MPORT_216_en = reset;
  assign ram_0_MPORT_217_data = 2'h0;
  assign ram_0_MPORT_217_addr = 8'hd9;
  assign ram_0_MPORT_217_mask = 1'h1;
  assign ram_0_MPORT_217_en = reset;
  assign ram_0_MPORT_218_data = 2'h0;
  assign ram_0_MPORT_218_addr = 8'hda;
  assign ram_0_MPORT_218_mask = 1'h1;
  assign ram_0_MPORT_218_en = reset;
  assign ram_0_MPORT_219_data = 2'h0;
  assign ram_0_MPORT_219_addr = 8'hdb;
  assign ram_0_MPORT_219_mask = 1'h1;
  assign ram_0_MPORT_219_en = reset;
  assign ram_0_MPORT_220_data = 2'h0;
  assign ram_0_MPORT_220_addr = 8'hdc;
  assign ram_0_MPORT_220_mask = 1'h1;
  assign ram_0_MPORT_220_en = reset;
  assign ram_0_MPORT_221_data = 2'h0;
  assign ram_0_MPORT_221_addr = 8'hdd;
  assign ram_0_MPORT_221_mask = 1'h1;
  assign ram_0_MPORT_221_en = reset;
  assign ram_0_MPORT_222_data = 2'h0;
  assign ram_0_MPORT_222_addr = 8'hde;
  assign ram_0_MPORT_222_mask = 1'h1;
  assign ram_0_MPORT_222_en = reset;
  assign ram_0_MPORT_223_data = 2'h0;
  assign ram_0_MPORT_223_addr = 8'hdf;
  assign ram_0_MPORT_223_mask = 1'h1;
  assign ram_0_MPORT_223_en = reset;
  assign ram_0_MPORT_224_data = 2'h0;
  assign ram_0_MPORT_224_addr = 8'he0;
  assign ram_0_MPORT_224_mask = 1'h1;
  assign ram_0_MPORT_224_en = reset;
  assign ram_0_MPORT_225_data = 2'h0;
  assign ram_0_MPORT_225_addr = 8'he1;
  assign ram_0_MPORT_225_mask = 1'h1;
  assign ram_0_MPORT_225_en = reset;
  assign ram_0_MPORT_226_data = 2'h0;
  assign ram_0_MPORT_226_addr = 8'he2;
  assign ram_0_MPORT_226_mask = 1'h1;
  assign ram_0_MPORT_226_en = reset;
  assign ram_0_MPORT_227_data = 2'h0;
  assign ram_0_MPORT_227_addr = 8'he3;
  assign ram_0_MPORT_227_mask = 1'h1;
  assign ram_0_MPORT_227_en = reset;
  assign ram_0_MPORT_228_data = 2'h0;
  assign ram_0_MPORT_228_addr = 8'he4;
  assign ram_0_MPORT_228_mask = 1'h1;
  assign ram_0_MPORT_228_en = reset;
  assign ram_0_MPORT_229_data = 2'h0;
  assign ram_0_MPORT_229_addr = 8'he5;
  assign ram_0_MPORT_229_mask = 1'h1;
  assign ram_0_MPORT_229_en = reset;
  assign ram_0_MPORT_230_data = 2'h0;
  assign ram_0_MPORT_230_addr = 8'he6;
  assign ram_0_MPORT_230_mask = 1'h1;
  assign ram_0_MPORT_230_en = reset;
  assign ram_0_MPORT_231_data = 2'h0;
  assign ram_0_MPORT_231_addr = 8'he7;
  assign ram_0_MPORT_231_mask = 1'h1;
  assign ram_0_MPORT_231_en = reset;
  assign ram_0_MPORT_232_data = 2'h0;
  assign ram_0_MPORT_232_addr = 8'he8;
  assign ram_0_MPORT_232_mask = 1'h1;
  assign ram_0_MPORT_232_en = reset;
  assign ram_0_MPORT_233_data = 2'h0;
  assign ram_0_MPORT_233_addr = 8'he9;
  assign ram_0_MPORT_233_mask = 1'h1;
  assign ram_0_MPORT_233_en = reset;
  assign ram_0_MPORT_234_data = 2'h0;
  assign ram_0_MPORT_234_addr = 8'hea;
  assign ram_0_MPORT_234_mask = 1'h1;
  assign ram_0_MPORT_234_en = reset;
  assign ram_0_MPORT_235_data = 2'h0;
  assign ram_0_MPORT_235_addr = 8'heb;
  assign ram_0_MPORT_235_mask = 1'h1;
  assign ram_0_MPORT_235_en = reset;
  assign ram_0_MPORT_236_data = 2'h0;
  assign ram_0_MPORT_236_addr = 8'hec;
  assign ram_0_MPORT_236_mask = 1'h1;
  assign ram_0_MPORT_236_en = reset;
  assign ram_0_MPORT_237_data = 2'h0;
  assign ram_0_MPORT_237_addr = 8'hed;
  assign ram_0_MPORT_237_mask = 1'h1;
  assign ram_0_MPORT_237_en = reset;
  assign ram_0_MPORT_238_data = 2'h0;
  assign ram_0_MPORT_238_addr = 8'hee;
  assign ram_0_MPORT_238_mask = 1'h1;
  assign ram_0_MPORT_238_en = reset;
  assign ram_0_MPORT_239_data = 2'h0;
  assign ram_0_MPORT_239_addr = 8'hef;
  assign ram_0_MPORT_239_mask = 1'h1;
  assign ram_0_MPORT_239_en = reset;
  assign ram_0_MPORT_240_data = 2'h0;
  assign ram_0_MPORT_240_addr = 8'hf0;
  assign ram_0_MPORT_240_mask = 1'h1;
  assign ram_0_MPORT_240_en = reset;
  assign ram_0_MPORT_241_data = 2'h0;
  assign ram_0_MPORT_241_addr = 8'hf1;
  assign ram_0_MPORT_241_mask = 1'h1;
  assign ram_0_MPORT_241_en = reset;
  assign ram_0_MPORT_242_data = 2'h0;
  assign ram_0_MPORT_242_addr = 8'hf2;
  assign ram_0_MPORT_242_mask = 1'h1;
  assign ram_0_MPORT_242_en = reset;
  assign ram_0_MPORT_243_data = 2'h0;
  assign ram_0_MPORT_243_addr = 8'hf3;
  assign ram_0_MPORT_243_mask = 1'h1;
  assign ram_0_MPORT_243_en = reset;
  assign ram_0_MPORT_244_data = 2'h0;
  assign ram_0_MPORT_244_addr = 8'hf4;
  assign ram_0_MPORT_244_mask = 1'h1;
  assign ram_0_MPORT_244_en = reset;
  assign ram_0_MPORT_245_data = 2'h0;
  assign ram_0_MPORT_245_addr = 8'hf5;
  assign ram_0_MPORT_245_mask = 1'h1;
  assign ram_0_MPORT_245_en = reset;
  assign ram_0_MPORT_246_data = 2'h0;
  assign ram_0_MPORT_246_addr = 8'hf6;
  assign ram_0_MPORT_246_mask = 1'h1;
  assign ram_0_MPORT_246_en = reset;
  assign ram_0_MPORT_247_data = 2'h0;
  assign ram_0_MPORT_247_addr = 8'hf7;
  assign ram_0_MPORT_247_mask = 1'h1;
  assign ram_0_MPORT_247_en = reset;
  assign ram_0_MPORT_248_data = 2'h0;
  assign ram_0_MPORT_248_addr = 8'hf8;
  assign ram_0_MPORT_248_mask = 1'h1;
  assign ram_0_MPORT_248_en = reset;
  assign ram_0_MPORT_249_data = 2'h0;
  assign ram_0_MPORT_249_addr = 8'hf9;
  assign ram_0_MPORT_249_mask = 1'h1;
  assign ram_0_MPORT_249_en = reset;
  assign ram_0_MPORT_250_data = 2'h0;
  assign ram_0_MPORT_250_addr = 8'hfa;
  assign ram_0_MPORT_250_mask = 1'h1;
  assign ram_0_MPORT_250_en = reset;
  assign ram_0_MPORT_251_data = 2'h0;
  assign ram_0_MPORT_251_addr = 8'hfb;
  assign ram_0_MPORT_251_mask = 1'h1;
  assign ram_0_MPORT_251_en = reset;
  assign ram_0_MPORT_252_data = 2'h0;
  assign ram_0_MPORT_252_addr = 8'hfc;
  assign ram_0_MPORT_252_mask = 1'h1;
  assign ram_0_MPORT_252_en = reset;
  assign ram_0_MPORT_253_data = 2'h0;
  assign ram_0_MPORT_253_addr = 8'hfd;
  assign ram_0_MPORT_253_mask = 1'h1;
  assign ram_0_MPORT_253_en = reset;
  assign ram_0_MPORT_254_data = 2'h0;
  assign ram_0_MPORT_254_addr = 8'hfe;
  assign ram_0_MPORT_254_mask = 1'h1;
  assign ram_0_MPORT_254_en = reset;
  assign ram_0_MPORT_255_data = 2'h0;
  assign ram_0_MPORT_255_addr = 8'hff;
  assign ram_0_MPORT_255_mask = 1'h1;
  assign ram_0_MPORT_255_en = reset;
  assign ram_0_MPORT_256_data = io_wdata[1:0];
  assign ram_0_MPORT_256_addr = io_addr;
  assign ram_0_MPORT_256_mask = io_wmask[0];
  assign ram_0_MPORT_256_en = io_rw;
  assign ram_1_io_rdata_MPORT_en = ram_1_io_rdata_MPORT_en_pipe_0;
  assign ram_1_io_rdata_MPORT_addr = ram_1_io_rdata_MPORT_addr_pipe_0;
  assign ram_1_io_rdata_MPORT_data = ram_1[ram_1_io_rdata_MPORT_addr]; // @[SRAM.scala 36:26]
  assign ram_1_MPORT_data = 2'h0;
  assign ram_1_MPORT_addr = 8'h0;
  assign ram_1_MPORT_mask = 1'h1;
  assign ram_1_MPORT_en = reset;
  assign ram_1_MPORT_1_data = 2'h0;
  assign ram_1_MPORT_1_addr = 8'h1;
  assign ram_1_MPORT_1_mask = 1'h1;
  assign ram_1_MPORT_1_en = reset;
  assign ram_1_MPORT_2_data = 2'h0;
  assign ram_1_MPORT_2_addr = 8'h2;
  assign ram_1_MPORT_2_mask = 1'h1;
  assign ram_1_MPORT_2_en = reset;
  assign ram_1_MPORT_3_data = 2'h0;
  assign ram_1_MPORT_3_addr = 8'h3;
  assign ram_1_MPORT_3_mask = 1'h1;
  assign ram_1_MPORT_3_en = reset;
  assign ram_1_MPORT_4_data = 2'h0;
  assign ram_1_MPORT_4_addr = 8'h4;
  assign ram_1_MPORT_4_mask = 1'h1;
  assign ram_1_MPORT_4_en = reset;
  assign ram_1_MPORT_5_data = 2'h0;
  assign ram_1_MPORT_5_addr = 8'h5;
  assign ram_1_MPORT_5_mask = 1'h1;
  assign ram_1_MPORT_5_en = reset;
  assign ram_1_MPORT_6_data = 2'h0;
  assign ram_1_MPORT_6_addr = 8'h6;
  assign ram_1_MPORT_6_mask = 1'h1;
  assign ram_1_MPORT_6_en = reset;
  assign ram_1_MPORT_7_data = 2'h0;
  assign ram_1_MPORT_7_addr = 8'h7;
  assign ram_1_MPORT_7_mask = 1'h1;
  assign ram_1_MPORT_7_en = reset;
  assign ram_1_MPORT_8_data = 2'h0;
  assign ram_1_MPORT_8_addr = 8'h8;
  assign ram_1_MPORT_8_mask = 1'h1;
  assign ram_1_MPORT_8_en = reset;
  assign ram_1_MPORT_9_data = 2'h0;
  assign ram_1_MPORT_9_addr = 8'h9;
  assign ram_1_MPORT_9_mask = 1'h1;
  assign ram_1_MPORT_9_en = reset;
  assign ram_1_MPORT_10_data = 2'h0;
  assign ram_1_MPORT_10_addr = 8'ha;
  assign ram_1_MPORT_10_mask = 1'h1;
  assign ram_1_MPORT_10_en = reset;
  assign ram_1_MPORT_11_data = 2'h0;
  assign ram_1_MPORT_11_addr = 8'hb;
  assign ram_1_MPORT_11_mask = 1'h1;
  assign ram_1_MPORT_11_en = reset;
  assign ram_1_MPORT_12_data = 2'h0;
  assign ram_1_MPORT_12_addr = 8'hc;
  assign ram_1_MPORT_12_mask = 1'h1;
  assign ram_1_MPORT_12_en = reset;
  assign ram_1_MPORT_13_data = 2'h0;
  assign ram_1_MPORT_13_addr = 8'hd;
  assign ram_1_MPORT_13_mask = 1'h1;
  assign ram_1_MPORT_13_en = reset;
  assign ram_1_MPORT_14_data = 2'h0;
  assign ram_1_MPORT_14_addr = 8'he;
  assign ram_1_MPORT_14_mask = 1'h1;
  assign ram_1_MPORT_14_en = reset;
  assign ram_1_MPORT_15_data = 2'h0;
  assign ram_1_MPORT_15_addr = 8'hf;
  assign ram_1_MPORT_15_mask = 1'h1;
  assign ram_1_MPORT_15_en = reset;
  assign ram_1_MPORT_16_data = 2'h0;
  assign ram_1_MPORT_16_addr = 8'h10;
  assign ram_1_MPORT_16_mask = 1'h1;
  assign ram_1_MPORT_16_en = reset;
  assign ram_1_MPORT_17_data = 2'h0;
  assign ram_1_MPORT_17_addr = 8'h11;
  assign ram_1_MPORT_17_mask = 1'h1;
  assign ram_1_MPORT_17_en = reset;
  assign ram_1_MPORT_18_data = 2'h0;
  assign ram_1_MPORT_18_addr = 8'h12;
  assign ram_1_MPORT_18_mask = 1'h1;
  assign ram_1_MPORT_18_en = reset;
  assign ram_1_MPORT_19_data = 2'h0;
  assign ram_1_MPORT_19_addr = 8'h13;
  assign ram_1_MPORT_19_mask = 1'h1;
  assign ram_1_MPORT_19_en = reset;
  assign ram_1_MPORT_20_data = 2'h0;
  assign ram_1_MPORT_20_addr = 8'h14;
  assign ram_1_MPORT_20_mask = 1'h1;
  assign ram_1_MPORT_20_en = reset;
  assign ram_1_MPORT_21_data = 2'h0;
  assign ram_1_MPORT_21_addr = 8'h15;
  assign ram_1_MPORT_21_mask = 1'h1;
  assign ram_1_MPORT_21_en = reset;
  assign ram_1_MPORT_22_data = 2'h0;
  assign ram_1_MPORT_22_addr = 8'h16;
  assign ram_1_MPORT_22_mask = 1'h1;
  assign ram_1_MPORT_22_en = reset;
  assign ram_1_MPORT_23_data = 2'h0;
  assign ram_1_MPORT_23_addr = 8'h17;
  assign ram_1_MPORT_23_mask = 1'h1;
  assign ram_1_MPORT_23_en = reset;
  assign ram_1_MPORT_24_data = 2'h0;
  assign ram_1_MPORT_24_addr = 8'h18;
  assign ram_1_MPORT_24_mask = 1'h1;
  assign ram_1_MPORT_24_en = reset;
  assign ram_1_MPORT_25_data = 2'h0;
  assign ram_1_MPORT_25_addr = 8'h19;
  assign ram_1_MPORT_25_mask = 1'h1;
  assign ram_1_MPORT_25_en = reset;
  assign ram_1_MPORT_26_data = 2'h0;
  assign ram_1_MPORT_26_addr = 8'h1a;
  assign ram_1_MPORT_26_mask = 1'h1;
  assign ram_1_MPORT_26_en = reset;
  assign ram_1_MPORT_27_data = 2'h0;
  assign ram_1_MPORT_27_addr = 8'h1b;
  assign ram_1_MPORT_27_mask = 1'h1;
  assign ram_1_MPORT_27_en = reset;
  assign ram_1_MPORT_28_data = 2'h0;
  assign ram_1_MPORT_28_addr = 8'h1c;
  assign ram_1_MPORT_28_mask = 1'h1;
  assign ram_1_MPORT_28_en = reset;
  assign ram_1_MPORT_29_data = 2'h0;
  assign ram_1_MPORT_29_addr = 8'h1d;
  assign ram_1_MPORT_29_mask = 1'h1;
  assign ram_1_MPORT_29_en = reset;
  assign ram_1_MPORT_30_data = 2'h0;
  assign ram_1_MPORT_30_addr = 8'h1e;
  assign ram_1_MPORT_30_mask = 1'h1;
  assign ram_1_MPORT_30_en = reset;
  assign ram_1_MPORT_31_data = 2'h0;
  assign ram_1_MPORT_31_addr = 8'h1f;
  assign ram_1_MPORT_31_mask = 1'h1;
  assign ram_1_MPORT_31_en = reset;
  assign ram_1_MPORT_32_data = 2'h0;
  assign ram_1_MPORT_32_addr = 8'h20;
  assign ram_1_MPORT_32_mask = 1'h1;
  assign ram_1_MPORT_32_en = reset;
  assign ram_1_MPORT_33_data = 2'h0;
  assign ram_1_MPORT_33_addr = 8'h21;
  assign ram_1_MPORT_33_mask = 1'h1;
  assign ram_1_MPORT_33_en = reset;
  assign ram_1_MPORT_34_data = 2'h0;
  assign ram_1_MPORT_34_addr = 8'h22;
  assign ram_1_MPORT_34_mask = 1'h1;
  assign ram_1_MPORT_34_en = reset;
  assign ram_1_MPORT_35_data = 2'h0;
  assign ram_1_MPORT_35_addr = 8'h23;
  assign ram_1_MPORT_35_mask = 1'h1;
  assign ram_1_MPORT_35_en = reset;
  assign ram_1_MPORT_36_data = 2'h0;
  assign ram_1_MPORT_36_addr = 8'h24;
  assign ram_1_MPORT_36_mask = 1'h1;
  assign ram_1_MPORT_36_en = reset;
  assign ram_1_MPORT_37_data = 2'h0;
  assign ram_1_MPORT_37_addr = 8'h25;
  assign ram_1_MPORT_37_mask = 1'h1;
  assign ram_1_MPORT_37_en = reset;
  assign ram_1_MPORT_38_data = 2'h0;
  assign ram_1_MPORT_38_addr = 8'h26;
  assign ram_1_MPORT_38_mask = 1'h1;
  assign ram_1_MPORT_38_en = reset;
  assign ram_1_MPORT_39_data = 2'h0;
  assign ram_1_MPORT_39_addr = 8'h27;
  assign ram_1_MPORT_39_mask = 1'h1;
  assign ram_1_MPORT_39_en = reset;
  assign ram_1_MPORT_40_data = 2'h0;
  assign ram_1_MPORT_40_addr = 8'h28;
  assign ram_1_MPORT_40_mask = 1'h1;
  assign ram_1_MPORT_40_en = reset;
  assign ram_1_MPORT_41_data = 2'h0;
  assign ram_1_MPORT_41_addr = 8'h29;
  assign ram_1_MPORT_41_mask = 1'h1;
  assign ram_1_MPORT_41_en = reset;
  assign ram_1_MPORT_42_data = 2'h0;
  assign ram_1_MPORT_42_addr = 8'h2a;
  assign ram_1_MPORT_42_mask = 1'h1;
  assign ram_1_MPORT_42_en = reset;
  assign ram_1_MPORT_43_data = 2'h0;
  assign ram_1_MPORT_43_addr = 8'h2b;
  assign ram_1_MPORT_43_mask = 1'h1;
  assign ram_1_MPORT_43_en = reset;
  assign ram_1_MPORT_44_data = 2'h0;
  assign ram_1_MPORT_44_addr = 8'h2c;
  assign ram_1_MPORT_44_mask = 1'h1;
  assign ram_1_MPORT_44_en = reset;
  assign ram_1_MPORT_45_data = 2'h0;
  assign ram_1_MPORT_45_addr = 8'h2d;
  assign ram_1_MPORT_45_mask = 1'h1;
  assign ram_1_MPORT_45_en = reset;
  assign ram_1_MPORT_46_data = 2'h0;
  assign ram_1_MPORT_46_addr = 8'h2e;
  assign ram_1_MPORT_46_mask = 1'h1;
  assign ram_1_MPORT_46_en = reset;
  assign ram_1_MPORT_47_data = 2'h0;
  assign ram_1_MPORT_47_addr = 8'h2f;
  assign ram_1_MPORT_47_mask = 1'h1;
  assign ram_1_MPORT_47_en = reset;
  assign ram_1_MPORT_48_data = 2'h0;
  assign ram_1_MPORT_48_addr = 8'h30;
  assign ram_1_MPORT_48_mask = 1'h1;
  assign ram_1_MPORT_48_en = reset;
  assign ram_1_MPORT_49_data = 2'h0;
  assign ram_1_MPORT_49_addr = 8'h31;
  assign ram_1_MPORT_49_mask = 1'h1;
  assign ram_1_MPORT_49_en = reset;
  assign ram_1_MPORT_50_data = 2'h0;
  assign ram_1_MPORT_50_addr = 8'h32;
  assign ram_1_MPORT_50_mask = 1'h1;
  assign ram_1_MPORT_50_en = reset;
  assign ram_1_MPORT_51_data = 2'h0;
  assign ram_1_MPORT_51_addr = 8'h33;
  assign ram_1_MPORT_51_mask = 1'h1;
  assign ram_1_MPORT_51_en = reset;
  assign ram_1_MPORT_52_data = 2'h0;
  assign ram_1_MPORT_52_addr = 8'h34;
  assign ram_1_MPORT_52_mask = 1'h1;
  assign ram_1_MPORT_52_en = reset;
  assign ram_1_MPORT_53_data = 2'h0;
  assign ram_1_MPORT_53_addr = 8'h35;
  assign ram_1_MPORT_53_mask = 1'h1;
  assign ram_1_MPORT_53_en = reset;
  assign ram_1_MPORT_54_data = 2'h0;
  assign ram_1_MPORT_54_addr = 8'h36;
  assign ram_1_MPORT_54_mask = 1'h1;
  assign ram_1_MPORT_54_en = reset;
  assign ram_1_MPORT_55_data = 2'h0;
  assign ram_1_MPORT_55_addr = 8'h37;
  assign ram_1_MPORT_55_mask = 1'h1;
  assign ram_1_MPORT_55_en = reset;
  assign ram_1_MPORT_56_data = 2'h0;
  assign ram_1_MPORT_56_addr = 8'h38;
  assign ram_1_MPORT_56_mask = 1'h1;
  assign ram_1_MPORT_56_en = reset;
  assign ram_1_MPORT_57_data = 2'h0;
  assign ram_1_MPORT_57_addr = 8'h39;
  assign ram_1_MPORT_57_mask = 1'h1;
  assign ram_1_MPORT_57_en = reset;
  assign ram_1_MPORT_58_data = 2'h0;
  assign ram_1_MPORT_58_addr = 8'h3a;
  assign ram_1_MPORT_58_mask = 1'h1;
  assign ram_1_MPORT_58_en = reset;
  assign ram_1_MPORT_59_data = 2'h0;
  assign ram_1_MPORT_59_addr = 8'h3b;
  assign ram_1_MPORT_59_mask = 1'h1;
  assign ram_1_MPORT_59_en = reset;
  assign ram_1_MPORT_60_data = 2'h0;
  assign ram_1_MPORT_60_addr = 8'h3c;
  assign ram_1_MPORT_60_mask = 1'h1;
  assign ram_1_MPORT_60_en = reset;
  assign ram_1_MPORT_61_data = 2'h0;
  assign ram_1_MPORT_61_addr = 8'h3d;
  assign ram_1_MPORT_61_mask = 1'h1;
  assign ram_1_MPORT_61_en = reset;
  assign ram_1_MPORT_62_data = 2'h0;
  assign ram_1_MPORT_62_addr = 8'h3e;
  assign ram_1_MPORT_62_mask = 1'h1;
  assign ram_1_MPORT_62_en = reset;
  assign ram_1_MPORT_63_data = 2'h0;
  assign ram_1_MPORT_63_addr = 8'h3f;
  assign ram_1_MPORT_63_mask = 1'h1;
  assign ram_1_MPORT_63_en = reset;
  assign ram_1_MPORT_64_data = 2'h0;
  assign ram_1_MPORT_64_addr = 8'h40;
  assign ram_1_MPORT_64_mask = 1'h1;
  assign ram_1_MPORT_64_en = reset;
  assign ram_1_MPORT_65_data = 2'h0;
  assign ram_1_MPORT_65_addr = 8'h41;
  assign ram_1_MPORT_65_mask = 1'h1;
  assign ram_1_MPORT_65_en = reset;
  assign ram_1_MPORT_66_data = 2'h0;
  assign ram_1_MPORT_66_addr = 8'h42;
  assign ram_1_MPORT_66_mask = 1'h1;
  assign ram_1_MPORT_66_en = reset;
  assign ram_1_MPORT_67_data = 2'h0;
  assign ram_1_MPORT_67_addr = 8'h43;
  assign ram_1_MPORT_67_mask = 1'h1;
  assign ram_1_MPORT_67_en = reset;
  assign ram_1_MPORT_68_data = 2'h0;
  assign ram_1_MPORT_68_addr = 8'h44;
  assign ram_1_MPORT_68_mask = 1'h1;
  assign ram_1_MPORT_68_en = reset;
  assign ram_1_MPORT_69_data = 2'h0;
  assign ram_1_MPORT_69_addr = 8'h45;
  assign ram_1_MPORT_69_mask = 1'h1;
  assign ram_1_MPORT_69_en = reset;
  assign ram_1_MPORT_70_data = 2'h0;
  assign ram_1_MPORT_70_addr = 8'h46;
  assign ram_1_MPORT_70_mask = 1'h1;
  assign ram_1_MPORT_70_en = reset;
  assign ram_1_MPORT_71_data = 2'h0;
  assign ram_1_MPORT_71_addr = 8'h47;
  assign ram_1_MPORT_71_mask = 1'h1;
  assign ram_1_MPORT_71_en = reset;
  assign ram_1_MPORT_72_data = 2'h0;
  assign ram_1_MPORT_72_addr = 8'h48;
  assign ram_1_MPORT_72_mask = 1'h1;
  assign ram_1_MPORT_72_en = reset;
  assign ram_1_MPORT_73_data = 2'h0;
  assign ram_1_MPORT_73_addr = 8'h49;
  assign ram_1_MPORT_73_mask = 1'h1;
  assign ram_1_MPORT_73_en = reset;
  assign ram_1_MPORT_74_data = 2'h0;
  assign ram_1_MPORT_74_addr = 8'h4a;
  assign ram_1_MPORT_74_mask = 1'h1;
  assign ram_1_MPORT_74_en = reset;
  assign ram_1_MPORT_75_data = 2'h0;
  assign ram_1_MPORT_75_addr = 8'h4b;
  assign ram_1_MPORT_75_mask = 1'h1;
  assign ram_1_MPORT_75_en = reset;
  assign ram_1_MPORT_76_data = 2'h0;
  assign ram_1_MPORT_76_addr = 8'h4c;
  assign ram_1_MPORT_76_mask = 1'h1;
  assign ram_1_MPORT_76_en = reset;
  assign ram_1_MPORT_77_data = 2'h0;
  assign ram_1_MPORT_77_addr = 8'h4d;
  assign ram_1_MPORT_77_mask = 1'h1;
  assign ram_1_MPORT_77_en = reset;
  assign ram_1_MPORT_78_data = 2'h0;
  assign ram_1_MPORT_78_addr = 8'h4e;
  assign ram_1_MPORT_78_mask = 1'h1;
  assign ram_1_MPORT_78_en = reset;
  assign ram_1_MPORT_79_data = 2'h0;
  assign ram_1_MPORT_79_addr = 8'h4f;
  assign ram_1_MPORT_79_mask = 1'h1;
  assign ram_1_MPORT_79_en = reset;
  assign ram_1_MPORT_80_data = 2'h0;
  assign ram_1_MPORT_80_addr = 8'h50;
  assign ram_1_MPORT_80_mask = 1'h1;
  assign ram_1_MPORT_80_en = reset;
  assign ram_1_MPORT_81_data = 2'h0;
  assign ram_1_MPORT_81_addr = 8'h51;
  assign ram_1_MPORT_81_mask = 1'h1;
  assign ram_1_MPORT_81_en = reset;
  assign ram_1_MPORT_82_data = 2'h0;
  assign ram_1_MPORT_82_addr = 8'h52;
  assign ram_1_MPORT_82_mask = 1'h1;
  assign ram_1_MPORT_82_en = reset;
  assign ram_1_MPORT_83_data = 2'h0;
  assign ram_1_MPORT_83_addr = 8'h53;
  assign ram_1_MPORT_83_mask = 1'h1;
  assign ram_1_MPORT_83_en = reset;
  assign ram_1_MPORT_84_data = 2'h0;
  assign ram_1_MPORT_84_addr = 8'h54;
  assign ram_1_MPORT_84_mask = 1'h1;
  assign ram_1_MPORT_84_en = reset;
  assign ram_1_MPORT_85_data = 2'h0;
  assign ram_1_MPORT_85_addr = 8'h55;
  assign ram_1_MPORT_85_mask = 1'h1;
  assign ram_1_MPORT_85_en = reset;
  assign ram_1_MPORT_86_data = 2'h0;
  assign ram_1_MPORT_86_addr = 8'h56;
  assign ram_1_MPORT_86_mask = 1'h1;
  assign ram_1_MPORT_86_en = reset;
  assign ram_1_MPORT_87_data = 2'h0;
  assign ram_1_MPORT_87_addr = 8'h57;
  assign ram_1_MPORT_87_mask = 1'h1;
  assign ram_1_MPORT_87_en = reset;
  assign ram_1_MPORT_88_data = 2'h0;
  assign ram_1_MPORT_88_addr = 8'h58;
  assign ram_1_MPORT_88_mask = 1'h1;
  assign ram_1_MPORT_88_en = reset;
  assign ram_1_MPORT_89_data = 2'h0;
  assign ram_1_MPORT_89_addr = 8'h59;
  assign ram_1_MPORT_89_mask = 1'h1;
  assign ram_1_MPORT_89_en = reset;
  assign ram_1_MPORT_90_data = 2'h0;
  assign ram_1_MPORT_90_addr = 8'h5a;
  assign ram_1_MPORT_90_mask = 1'h1;
  assign ram_1_MPORT_90_en = reset;
  assign ram_1_MPORT_91_data = 2'h0;
  assign ram_1_MPORT_91_addr = 8'h5b;
  assign ram_1_MPORT_91_mask = 1'h1;
  assign ram_1_MPORT_91_en = reset;
  assign ram_1_MPORT_92_data = 2'h0;
  assign ram_1_MPORT_92_addr = 8'h5c;
  assign ram_1_MPORT_92_mask = 1'h1;
  assign ram_1_MPORT_92_en = reset;
  assign ram_1_MPORT_93_data = 2'h0;
  assign ram_1_MPORT_93_addr = 8'h5d;
  assign ram_1_MPORT_93_mask = 1'h1;
  assign ram_1_MPORT_93_en = reset;
  assign ram_1_MPORT_94_data = 2'h0;
  assign ram_1_MPORT_94_addr = 8'h5e;
  assign ram_1_MPORT_94_mask = 1'h1;
  assign ram_1_MPORT_94_en = reset;
  assign ram_1_MPORT_95_data = 2'h0;
  assign ram_1_MPORT_95_addr = 8'h5f;
  assign ram_1_MPORT_95_mask = 1'h1;
  assign ram_1_MPORT_95_en = reset;
  assign ram_1_MPORT_96_data = 2'h0;
  assign ram_1_MPORT_96_addr = 8'h60;
  assign ram_1_MPORT_96_mask = 1'h1;
  assign ram_1_MPORT_96_en = reset;
  assign ram_1_MPORT_97_data = 2'h0;
  assign ram_1_MPORT_97_addr = 8'h61;
  assign ram_1_MPORT_97_mask = 1'h1;
  assign ram_1_MPORT_97_en = reset;
  assign ram_1_MPORT_98_data = 2'h0;
  assign ram_1_MPORT_98_addr = 8'h62;
  assign ram_1_MPORT_98_mask = 1'h1;
  assign ram_1_MPORT_98_en = reset;
  assign ram_1_MPORT_99_data = 2'h0;
  assign ram_1_MPORT_99_addr = 8'h63;
  assign ram_1_MPORT_99_mask = 1'h1;
  assign ram_1_MPORT_99_en = reset;
  assign ram_1_MPORT_100_data = 2'h0;
  assign ram_1_MPORT_100_addr = 8'h64;
  assign ram_1_MPORT_100_mask = 1'h1;
  assign ram_1_MPORT_100_en = reset;
  assign ram_1_MPORT_101_data = 2'h0;
  assign ram_1_MPORT_101_addr = 8'h65;
  assign ram_1_MPORT_101_mask = 1'h1;
  assign ram_1_MPORT_101_en = reset;
  assign ram_1_MPORT_102_data = 2'h0;
  assign ram_1_MPORT_102_addr = 8'h66;
  assign ram_1_MPORT_102_mask = 1'h1;
  assign ram_1_MPORT_102_en = reset;
  assign ram_1_MPORT_103_data = 2'h0;
  assign ram_1_MPORT_103_addr = 8'h67;
  assign ram_1_MPORT_103_mask = 1'h1;
  assign ram_1_MPORT_103_en = reset;
  assign ram_1_MPORT_104_data = 2'h0;
  assign ram_1_MPORT_104_addr = 8'h68;
  assign ram_1_MPORT_104_mask = 1'h1;
  assign ram_1_MPORT_104_en = reset;
  assign ram_1_MPORT_105_data = 2'h0;
  assign ram_1_MPORT_105_addr = 8'h69;
  assign ram_1_MPORT_105_mask = 1'h1;
  assign ram_1_MPORT_105_en = reset;
  assign ram_1_MPORT_106_data = 2'h0;
  assign ram_1_MPORT_106_addr = 8'h6a;
  assign ram_1_MPORT_106_mask = 1'h1;
  assign ram_1_MPORT_106_en = reset;
  assign ram_1_MPORT_107_data = 2'h0;
  assign ram_1_MPORT_107_addr = 8'h6b;
  assign ram_1_MPORT_107_mask = 1'h1;
  assign ram_1_MPORT_107_en = reset;
  assign ram_1_MPORT_108_data = 2'h0;
  assign ram_1_MPORT_108_addr = 8'h6c;
  assign ram_1_MPORT_108_mask = 1'h1;
  assign ram_1_MPORT_108_en = reset;
  assign ram_1_MPORT_109_data = 2'h0;
  assign ram_1_MPORT_109_addr = 8'h6d;
  assign ram_1_MPORT_109_mask = 1'h1;
  assign ram_1_MPORT_109_en = reset;
  assign ram_1_MPORT_110_data = 2'h0;
  assign ram_1_MPORT_110_addr = 8'h6e;
  assign ram_1_MPORT_110_mask = 1'h1;
  assign ram_1_MPORT_110_en = reset;
  assign ram_1_MPORT_111_data = 2'h0;
  assign ram_1_MPORT_111_addr = 8'h6f;
  assign ram_1_MPORT_111_mask = 1'h1;
  assign ram_1_MPORT_111_en = reset;
  assign ram_1_MPORT_112_data = 2'h0;
  assign ram_1_MPORT_112_addr = 8'h70;
  assign ram_1_MPORT_112_mask = 1'h1;
  assign ram_1_MPORT_112_en = reset;
  assign ram_1_MPORT_113_data = 2'h0;
  assign ram_1_MPORT_113_addr = 8'h71;
  assign ram_1_MPORT_113_mask = 1'h1;
  assign ram_1_MPORT_113_en = reset;
  assign ram_1_MPORT_114_data = 2'h0;
  assign ram_1_MPORT_114_addr = 8'h72;
  assign ram_1_MPORT_114_mask = 1'h1;
  assign ram_1_MPORT_114_en = reset;
  assign ram_1_MPORT_115_data = 2'h0;
  assign ram_1_MPORT_115_addr = 8'h73;
  assign ram_1_MPORT_115_mask = 1'h1;
  assign ram_1_MPORT_115_en = reset;
  assign ram_1_MPORT_116_data = 2'h0;
  assign ram_1_MPORT_116_addr = 8'h74;
  assign ram_1_MPORT_116_mask = 1'h1;
  assign ram_1_MPORT_116_en = reset;
  assign ram_1_MPORT_117_data = 2'h0;
  assign ram_1_MPORT_117_addr = 8'h75;
  assign ram_1_MPORT_117_mask = 1'h1;
  assign ram_1_MPORT_117_en = reset;
  assign ram_1_MPORT_118_data = 2'h0;
  assign ram_1_MPORT_118_addr = 8'h76;
  assign ram_1_MPORT_118_mask = 1'h1;
  assign ram_1_MPORT_118_en = reset;
  assign ram_1_MPORT_119_data = 2'h0;
  assign ram_1_MPORT_119_addr = 8'h77;
  assign ram_1_MPORT_119_mask = 1'h1;
  assign ram_1_MPORT_119_en = reset;
  assign ram_1_MPORT_120_data = 2'h0;
  assign ram_1_MPORT_120_addr = 8'h78;
  assign ram_1_MPORT_120_mask = 1'h1;
  assign ram_1_MPORT_120_en = reset;
  assign ram_1_MPORT_121_data = 2'h0;
  assign ram_1_MPORT_121_addr = 8'h79;
  assign ram_1_MPORT_121_mask = 1'h1;
  assign ram_1_MPORT_121_en = reset;
  assign ram_1_MPORT_122_data = 2'h0;
  assign ram_1_MPORT_122_addr = 8'h7a;
  assign ram_1_MPORT_122_mask = 1'h1;
  assign ram_1_MPORT_122_en = reset;
  assign ram_1_MPORT_123_data = 2'h0;
  assign ram_1_MPORT_123_addr = 8'h7b;
  assign ram_1_MPORT_123_mask = 1'h1;
  assign ram_1_MPORT_123_en = reset;
  assign ram_1_MPORT_124_data = 2'h0;
  assign ram_1_MPORT_124_addr = 8'h7c;
  assign ram_1_MPORT_124_mask = 1'h1;
  assign ram_1_MPORT_124_en = reset;
  assign ram_1_MPORT_125_data = 2'h0;
  assign ram_1_MPORT_125_addr = 8'h7d;
  assign ram_1_MPORT_125_mask = 1'h1;
  assign ram_1_MPORT_125_en = reset;
  assign ram_1_MPORT_126_data = 2'h0;
  assign ram_1_MPORT_126_addr = 8'h7e;
  assign ram_1_MPORT_126_mask = 1'h1;
  assign ram_1_MPORT_126_en = reset;
  assign ram_1_MPORT_127_data = 2'h0;
  assign ram_1_MPORT_127_addr = 8'h7f;
  assign ram_1_MPORT_127_mask = 1'h1;
  assign ram_1_MPORT_127_en = reset;
  assign ram_1_MPORT_128_data = 2'h0;
  assign ram_1_MPORT_128_addr = 8'h80;
  assign ram_1_MPORT_128_mask = 1'h1;
  assign ram_1_MPORT_128_en = reset;
  assign ram_1_MPORT_129_data = 2'h0;
  assign ram_1_MPORT_129_addr = 8'h81;
  assign ram_1_MPORT_129_mask = 1'h1;
  assign ram_1_MPORT_129_en = reset;
  assign ram_1_MPORT_130_data = 2'h0;
  assign ram_1_MPORT_130_addr = 8'h82;
  assign ram_1_MPORT_130_mask = 1'h1;
  assign ram_1_MPORT_130_en = reset;
  assign ram_1_MPORT_131_data = 2'h0;
  assign ram_1_MPORT_131_addr = 8'h83;
  assign ram_1_MPORT_131_mask = 1'h1;
  assign ram_1_MPORT_131_en = reset;
  assign ram_1_MPORT_132_data = 2'h0;
  assign ram_1_MPORT_132_addr = 8'h84;
  assign ram_1_MPORT_132_mask = 1'h1;
  assign ram_1_MPORT_132_en = reset;
  assign ram_1_MPORT_133_data = 2'h0;
  assign ram_1_MPORT_133_addr = 8'h85;
  assign ram_1_MPORT_133_mask = 1'h1;
  assign ram_1_MPORT_133_en = reset;
  assign ram_1_MPORT_134_data = 2'h0;
  assign ram_1_MPORT_134_addr = 8'h86;
  assign ram_1_MPORT_134_mask = 1'h1;
  assign ram_1_MPORT_134_en = reset;
  assign ram_1_MPORT_135_data = 2'h0;
  assign ram_1_MPORT_135_addr = 8'h87;
  assign ram_1_MPORT_135_mask = 1'h1;
  assign ram_1_MPORT_135_en = reset;
  assign ram_1_MPORT_136_data = 2'h0;
  assign ram_1_MPORT_136_addr = 8'h88;
  assign ram_1_MPORT_136_mask = 1'h1;
  assign ram_1_MPORT_136_en = reset;
  assign ram_1_MPORT_137_data = 2'h0;
  assign ram_1_MPORT_137_addr = 8'h89;
  assign ram_1_MPORT_137_mask = 1'h1;
  assign ram_1_MPORT_137_en = reset;
  assign ram_1_MPORT_138_data = 2'h0;
  assign ram_1_MPORT_138_addr = 8'h8a;
  assign ram_1_MPORT_138_mask = 1'h1;
  assign ram_1_MPORT_138_en = reset;
  assign ram_1_MPORT_139_data = 2'h0;
  assign ram_1_MPORT_139_addr = 8'h8b;
  assign ram_1_MPORT_139_mask = 1'h1;
  assign ram_1_MPORT_139_en = reset;
  assign ram_1_MPORT_140_data = 2'h0;
  assign ram_1_MPORT_140_addr = 8'h8c;
  assign ram_1_MPORT_140_mask = 1'h1;
  assign ram_1_MPORT_140_en = reset;
  assign ram_1_MPORT_141_data = 2'h0;
  assign ram_1_MPORT_141_addr = 8'h8d;
  assign ram_1_MPORT_141_mask = 1'h1;
  assign ram_1_MPORT_141_en = reset;
  assign ram_1_MPORT_142_data = 2'h0;
  assign ram_1_MPORT_142_addr = 8'h8e;
  assign ram_1_MPORT_142_mask = 1'h1;
  assign ram_1_MPORT_142_en = reset;
  assign ram_1_MPORT_143_data = 2'h0;
  assign ram_1_MPORT_143_addr = 8'h8f;
  assign ram_1_MPORT_143_mask = 1'h1;
  assign ram_1_MPORT_143_en = reset;
  assign ram_1_MPORT_144_data = 2'h0;
  assign ram_1_MPORT_144_addr = 8'h90;
  assign ram_1_MPORT_144_mask = 1'h1;
  assign ram_1_MPORT_144_en = reset;
  assign ram_1_MPORT_145_data = 2'h0;
  assign ram_1_MPORT_145_addr = 8'h91;
  assign ram_1_MPORT_145_mask = 1'h1;
  assign ram_1_MPORT_145_en = reset;
  assign ram_1_MPORT_146_data = 2'h0;
  assign ram_1_MPORT_146_addr = 8'h92;
  assign ram_1_MPORT_146_mask = 1'h1;
  assign ram_1_MPORT_146_en = reset;
  assign ram_1_MPORT_147_data = 2'h0;
  assign ram_1_MPORT_147_addr = 8'h93;
  assign ram_1_MPORT_147_mask = 1'h1;
  assign ram_1_MPORT_147_en = reset;
  assign ram_1_MPORT_148_data = 2'h0;
  assign ram_1_MPORT_148_addr = 8'h94;
  assign ram_1_MPORT_148_mask = 1'h1;
  assign ram_1_MPORT_148_en = reset;
  assign ram_1_MPORT_149_data = 2'h0;
  assign ram_1_MPORT_149_addr = 8'h95;
  assign ram_1_MPORT_149_mask = 1'h1;
  assign ram_1_MPORT_149_en = reset;
  assign ram_1_MPORT_150_data = 2'h0;
  assign ram_1_MPORT_150_addr = 8'h96;
  assign ram_1_MPORT_150_mask = 1'h1;
  assign ram_1_MPORT_150_en = reset;
  assign ram_1_MPORT_151_data = 2'h0;
  assign ram_1_MPORT_151_addr = 8'h97;
  assign ram_1_MPORT_151_mask = 1'h1;
  assign ram_1_MPORT_151_en = reset;
  assign ram_1_MPORT_152_data = 2'h0;
  assign ram_1_MPORT_152_addr = 8'h98;
  assign ram_1_MPORT_152_mask = 1'h1;
  assign ram_1_MPORT_152_en = reset;
  assign ram_1_MPORT_153_data = 2'h0;
  assign ram_1_MPORT_153_addr = 8'h99;
  assign ram_1_MPORT_153_mask = 1'h1;
  assign ram_1_MPORT_153_en = reset;
  assign ram_1_MPORT_154_data = 2'h0;
  assign ram_1_MPORT_154_addr = 8'h9a;
  assign ram_1_MPORT_154_mask = 1'h1;
  assign ram_1_MPORT_154_en = reset;
  assign ram_1_MPORT_155_data = 2'h0;
  assign ram_1_MPORT_155_addr = 8'h9b;
  assign ram_1_MPORT_155_mask = 1'h1;
  assign ram_1_MPORT_155_en = reset;
  assign ram_1_MPORT_156_data = 2'h0;
  assign ram_1_MPORT_156_addr = 8'h9c;
  assign ram_1_MPORT_156_mask = 1'h1;
  assign ram_1_MPORT_156_en = reset;
  assign ram_1_MPORT_157_data = 2'h0;
  assign ram_1_MPORT_157_addr = 8'h9d;
  assign ram_1_MPORT_157_mask = 1'h1;
  assign ram_1_MPORT_157_en = reset;
  assign ram_1_MPORT_158_data = 2'h0;
  assign ram_1_MPORT_158_addr = 8'h9e;
  assign ram_1_MPORT_158_mask = 1'h1;
  assign ram_1_MPORT_158_en = reset;
  assign ram_1_MPORT_159_data = 2'h0;
  assign ram_1_MPORT_159_addr = 8'h9f;
  assign ram_1_MPORT_159_mask = 1'h1;
  assign ram_1_MPORT_159_en = reset;
  assign ram_1_MPORT_160_data = 2'h0;
  assign ram_1_MPORT_160_addr = 8'ha0;
  assign ram_1_MPORT_160_mask = 1'h1;
  assign ram_1_MPORT_160_en = reset;
  assign ram_1_MPORT_161_data = 2'h0;
  assign ram_1_MPORT_161_addr = 8'ha1;
  assign ram_1_MPORT_161_mask = 1'h1;
  assign ram_1_MPORT_161_en = reset;
  assign ram_1_MPORT_162_data = 2'h0;
  assign ram_1_MPORT_162_addr = 8'ha2;
  assign ram_1_MPORT_162_mask = 1'h1;
  assign ram_1_MPORT_162_en = reset;
  assign ram_1_MPORT_163_data = 2'h0;
  assign ram_1_MPORT_163_addr = 8'ha3;
  assign ram_1_MPORT_163_mask = 1'h1;
  assign ram_1_MPORT_163_en = reset;
  assign ram_1_MPORT_164_data = 2'h0;
  assign ram_1_MPORT_164_addr = 8'ha4;
  assign ram_1_MPORT_164_mask = 1'h1;
  assign ram_1_MPORT_164_en = reset;
  assign ram_1_MPORT_165_data = 2'h0;
  assign ram_1_MPORT_165_addr = 8'ha5;
  assign ram_1_MPORT_165_mask = 1'h1;
  assign ram_1_MPORT_165_en = reset;
  assign ram_1_MPORT_166_data = 2'h0;
  assign ram_1_MPORT_166_addr = 8'ha6;
  assign ram_1_MPORT_166_mask = 1'h1;
  assign ram_1_MPORT_166_en = reset;
  assign ram_1_MPORT_167_data = 2'h0;
  assign ram_1_MPORT_167_addr = 8'ha7;
  assign ram_1_MPORT_167_mask = 1'h1;
  assign ram_1_MPORT_167_en = reset;
  assign ram_1_MPORT_168_data = 2'h0;
  assign ram_1_MPORT_168_addr = 8'ha8;
  assign ram_1_MPORT_168_mask = 1'h1;
  assign ram_1_MPORT_168_en = reset;
  assign ram_1_MPORT_169_data = 2'h0;
  assign ram_1_MPORT_169_addr = 8'ha9;
  assign ram_1_MPORT_169_mask = 1'h1;
  assign ram_1_MPORT_169_en = reset;
  assign ram_1_MPORT_170_data = 2'h0;
  assign ram_1_MPORT_170_addr = 8'haa;
  assign ram_1_MPORT_170_mask = 1'h1;
  assign ram_1_MPORT_170_en = reset;
  assign ram_1_MPORT_171_data = 2'h0;
  assign ram_1_MPORT_171_addr = 8'hab;
  assign ram_1_MPORT_171_mask = 1'h1;
  assign ram_1_MPORT_171_en = reset;
  assign ram_1_MPORT_172_data = 2'h0;
  assign ram_1_MPORT_172_addr = 8'hac;
  assign ram_1_MPORT_172_mask = 1'h1;
  assign ram_1_MPORT_172_en = reset;
  assign ram_1_MPORT_173_data = 2'h0;
  assign ram_1_MPORT_173_addr = 8'had;
  assign ram_1_MPORT_173_mask = 1'h1;
  assign ram_1_MPORT_173_en = reset;
  assign ram_1_MPORT_174_data = 2'h0;
  assign ram_1_MPORT_174_addr = 8'hae;
  assign ram_1_MPORT_174_mask = 1'h1;
  assign ram_1_MPORT_174_en = reset;
  assign ram_1_MPORT_175_data = 2'h0;
  assign ram_1_MPORT_175_addr = 8'haf;
  assign ram_1_MPORT_175_mask = 1'h1;
  assign ram_1_MPORT_175_en = reset;
  assign ram_1_MPORT_176_data = 2'h0;
  assign ram_1_MPORT_176_addr = 8'hb0;
  assign ram_1_MPORT_176_mask = 1'h1;
  assign ram_1_MPORT_176_en = reset;
  assign ram_1_MPORT_177_data = 2'h0;
  assign ram_1_MPORT_177_addr = 8'hb1;
  assign ram_1_MPORT_177_mask = 1'h1;
  assign ram_1_MPORT_177_en = reset;
  assign ram_1_MPORT_178_data = 2'h0;
  assign ram_1_MPORT_178_addr = 8'hb2;
  assign ram_1_MPORT_178_mask = 1'h1;
  assign ram_1_MPORT_178_en = reset;
  assign ram_1_MPORT_179_data = 2'h0;
  assign ram_1_MPORT_179_addr = 8'hb3;
  assign ram_1_MPORT_179_mask = 1'h1;
  assign ram_1_MPORT_179_en = reset;
  assign ram_1_MPORT_180_data = 2'h0;
  assign ram_1_MPORT_180_addr = 8'hb4;
  assign ram_1_MPORT_180_mask = 1'h1;
  assign ram_1_MPORT_180_en = reset;
  assign ram_1_MPORT_181_data = 2'h0;
  assign ram_1_MPORT_181_addr = 8'hb5;
  assign ram_1_MPORT_181_mask = 1'h1;
  assign ram_1_MPORT_181_en = reset;
  assign ram_1_MPORT_182_data = 2'h0;
  assign ram_1_MPORT_182_addr = 8'hb6;
  assign ram_1_MPORT_182_mask = 1'h1;
  assign ram_1_MPORT_182_en = reset;
  assign ram_1_MPORT_183_data = 2'h0;
  assign ram_1_MPORT_183_addr = 8'hb7;
  assign ram_1_MPORT_183_mask = 1'h1;
  assign ram_1_MPORT_183_en = reset;
  assign ram_1_MPORT_184_data = 2'h0;
  assign ram_1_MPORT_184_addr = 8'hb8;
  assign ram_1_MPORT_184_mask = 1'h1;
  assign ram_1_MPORT_184_en = reset;
  assign ram_1_MPORT_185_data = 2'h0;
  assign ram_1_MPORT_185_addr = 8'hb9;
  assign ram_1_MPORT_185_mask = 1'h1;
  assign ram_1_MPORT_185_en = reset;
  assign ram_1_MPORT_186_data = 2'h0;
  assign ram_1_MPORT_186_addr = 8'hba;
  assign ram_1_MPORT_186_mask = 1'h1;
  assign ram_1_MPORT_186_en = reset;
  assign ram_1_MPORT_187_data = 2'h0;
  assign ram_1_MPORT_187_addr = 8'hbb;
  assign ram_1_MPORT_187_mask = 1'h1;
  assign ram_1_MPORT_187_en = reset;
  assign ram_1_MPORT_188_data = 2'h0;
  assign ram_1_MPORT_188_addr = 8'hbc;
  assign ram_1_MPORT_188_mask = 1'h1;
  assign ram_1_MPORT_188_en = reset;
  assign ram_1_MPORT_189_data = 2'h0;
  assign ram_1_MPORT_189_addr = 8'hbd;
  assign ram_1_MPORT_189_mask = 1'h1;
  assign ram_1_MPORT_189_en = reset;
  assign ram_1_MPORT_190_data = 2'h0;
  assign ram_1_MPORT_190_addr = 8'hbe;
  assign ram_1_MPORT_190_mask = 1'h1;
  assign ram_1_MPORT_190_en = reset;
  assign ram_1_MPORT_191_data = 2'h0;
  assign ram_1_MPORT_191_addr = 8'hbf;
  assign ram_1_MPORT_191_mask = 1'h1;
  assign ram_1_MPORT_191_en = reset;
  assign ram_1_MPORT_192_data = 2'h0;
  assign ram_1_MPORT_192_addr = 8'hc0;
  assign ram_1_MPORT_192_mask = 1'h1;
  assign ram_1_MPORT_192_en = reset;
  assign ram_1_MPORT_193_data = 2'h0;
  assign ram_1_MPORT_193_addr = 8'hc1;
  assign ram_1_MPORT_193_mask = 1'h1;
  assign ram_1_MPORT_193_en = reset;
  assign ram_1_MPORT_194_data = 2'h0;
  assign ram_1_MPORT_194_addr = 8'hc2;
  assign ram_1_MPORT_194_mask = 1'h1;
  assign ram_1_MPORT_194_en = reset;
  assign ram_1_MPORT_195_data = 2'h0;
  assign ram_1_MPORT_195_addr = 8'hc3;
  assign ram_1_MPORT_195_mask = 1'h1;
  assign ram_1_MPORT_195_en = reset;
  assign ram_1_MPORT_196_data = 2'h0;
  assign ram_1_MPORT_196_addr = 8'hc4;
  assign ram_1_MPORT_196_mask = 1'h1;
  assign ram_1_MPORT_196_en = reset;
  assign ram_1_MPORT_197_data = 2'h0;
  assign ram_1_MPORT_197_addr = 8'hc5;
  assign ram_1_MPORT_197_mask = 1'h1;
  assign ram_1_MPORT_197_en = reset;
  assign ram_1_MPORT_198_data = 2'h0;
  assign ram_1_MPORT_198_addr = 8'hc6;
  assign ram_1_MPORT_198_mask = 1'h1;
  assign ram_1_MPORT_198_en = reset;
  assign ram_1_MPORT_199_data = 2'h0;
  assign ram_1_MPORT_199_addr = 8'hc7;
  assign ram_1_MPORT_199_mask = 1'h1;
  assign ram_1_MPORT_199_en = reset;
  assign ram_1_MPORT_200_data = 2'h0;
  assign ram_1_MPORT_200_addr = 8'hc8;
  assign ram_1_MPORT_200_mask = 1'h1;
  assign ram_1_MPORT_200_en = reset;
  assign ram_1_MPORT_201_data = 2'h0;
  assign ram_1_MPORT_201_addr = 8'hc9;
  assign ram_1_MPORT_201_mask = 1'h1;
  assign ram_1_MPORT_201_en = reset;
  assign ram_1_MPORT_202_data = 2'h0;
  assign ram_1_MPORT_202_addr = 8'hca;
  assign ram_1_MPORT_202_mask = 1'h1;
  assign ram_1_MPORT_202_en = reset;
  assign ram_1_MPORT_203_data = 2'h0;
  assign ram_1_MPORT_203_addr = 8'hcb;
  assign ram_1_MPORT_203_mask = 1'h1;
  assign ram_1_MPORT_203_en = reset;
  assign ram_1_MPORT_204_data = 2'h0;
  assign ram_1_MPORT_204_addr = 8'hcc;
  assign ram_1_MPORT_204_mask = 1'h1;
  assign ram_1_MPORT_204_en = reset;
  assign ram_1_MPORT_205_data = 2'h0;
  assign ram_1_MPORT_205_addr = 8'hcd;
  assign ram_1_MPORT_205_mask = 1'h1;
  assign ram_1_MPORT_205_en = reset;
  assign ram_1_MPORT_206_data = 2'h0;
  assign ram_1_MPORT_206_addr = 8'hce;
  assign ram_1_MPORT_206_mask = 1'h1;
  assign ram_1_MPORT_206_en = reset;
  assign ram_1_MPORT_207_data = 2'h0;
  assign ram_1_MPORT_207_addr = 8'hcf;
  assign ram_1_MPORT_207_mask = 1'h1;
  assign ram_1_MPORT_207_en = reset;
  assign ram_1_MPORT_208_data = 2'h0;
  assign ram_1_MPORT_208_addr = 8'hd0;
  assign ram_1_MPORT_208_mask = 1'h1;
  assign ram_1_MPORT_208_en = reset;
  assign ram_1_MPORT_209_data = 2'h0;
  assign ram_1_MPORT_209_addr = 8'hd1;
  assign ram_1_MPORT_209_mask = 1'h1;
  assign ram_1_MPORT_209_en = reset;
  assign ram_1_MPORT_210_data = 2'h0;
  assign ram_1_MPORT_210_addr = 8'hd2;
  assign ram_1_MPORT_210_mask = 1'h1;
  assign ram_1_MPORT_210_en = reset;
  assign ram_1_MPORT_211_data = 2'h0;
  assign ram_1_MPORT_211_addr = 8'hd3;
  assign ram_1_MPORT_211_mask = 1'h1;
  assign ram_1_MPORT_211_en = reset;
  assign ram_1_MPORT_212_data = 2'h0;
  assign ram_1_MPORT_212_addr = 8'hd4;
  assign ram_1_MPORT_212_mask = 1'h1;
  assign ram_1_MPORT_212_en = reset;
  assign ram_1_MPORT_213_data = 2'h0;
  assign ram_1_MPORT_213_addr = 8'hd5;
  assign ram_1_MPORT_213_mask = 1'h1;
  assign ram_1_MPORT_213_en = reset;
  assign ram_1_MPORT_214_data = 2'h0;
  assign ram_1_MPORT_214_addr = 8'hd6;
  assign ram_1_MPORT_214_mask = 1'h1;
  assign ram_1_MPORT_214_en = reset;
  assign ram_1_MPORT_215_data = 2'h0;
  assign ram_1_MPORT_215_addr = 8'hd7;
  assign ram_1_MPORT_215_mask = 1'h1;
  assign ram_1_MPORT_215_en = reset;
  assign ram_1_MPORT_216_data = 2'h0;
  assign ram_1_MPORT_216_addr = 8'hd8;
  assign ram_1_MPORT_216_mask = 1'h1;
  assign ram_1_MPORT_216_en = reset;
  assign ram_1_MPORT_217_data = 2'h0;
  assign ram_1_MPORT_217_addr = 8'hd9;
  assign ram_1_MPORT_217_mask = 1'h1;
  assign ram_1_MPORT_217_en = reset;
  assign ram_1_MPORT_218_data = 2'h0;
  assign ram_1_MPORT_218_addr = 8'hda;
  assign ram_1_MPORT_218_mask = 1'h1;
  assign ram_1_MPORT_218_en = reset;
  assign ram_1_MPORT_219_data = 2'h0;
  assign ram_1_MPORT_219_addr = 8'hdb;
  assign ram_1_MPORT_219_mask = 1'h1;
  assign ram_1_MPORT_219_en = reset;
  assign ram_1_MPORT_220_data = 2'h0;
  assign ram_1_MPORT_220_addr = 8'hdc;
  assign ram_1_MPORT_220_mask = 1'h1;
  assign ram_1_MPORT_220_en = reset;
  assign ram_1_MPORT_221_data = 2'h0;
  assign ram_1_MPORT_221_addr = 8'hdd;
  assign ram_1_MPORT_221_mask = 1'h1;
  assign ram_1_MPORT_221_en = reset;
  assign ram_1_MPORT_222_data = 2'h0;
  assign ram_1_MPORT_222_addr = 8'hde;
  assign ram_1_MPORT_222_mask = 1'h1;
  assign ram_1_MPORT_222_en = reset;
  assign ram_1_MPORT_223_data = 2'h0;
  assign ram_1_MPORT_223_addr = 8'hdf;
  assign ram_1_MPORT_223_mask = 1'h1;
  assign ram_1_MPORT_223_en = reset;
  assign ram_1_MPORT_224_data = 2'h0;
  assign ram_1_MPORT_224_addr = 8'he0;
  assign ram_1_MPORT_224_mask = 1'h1;
  assign ram_1_MPORT_224_en = reset;
  assign ram_1_MPORT_225_data = 2'h0;
  assign ram_1_MPORT_225_addr = 8'he1;
  assign ram_1_MPORT_225_mask = 1'h1;
  assign ram_1_MPORT_225_en = reset;
  assign ram_1_MPORT_226_data = 2'h0;
  assign ram_1_MPORT_226_addr = 8'he2;
  assign ram_1_MPORT_226_mask = 1'h1;
  assign ram_1_MPORT_226_en = reset;
  assign ram_1_MPORT_227_data = 2'h0;
  assign ram_1_MPORT_227_addr = 8'he3;
  assign ram_1_MPORT_227_mask = 1'h1;
  assign ram_1_MPORT_227_en = reset;
  assign ram_1_MPORT_228_data = 2'h0;
  assign ram_1_MPORT_228_addr = 8'he4;
  assign ram_1_MPORT_228_mask = 1'h1;
  assign ram_1_MPORT_228_en = reset;
  assign ram_1_MPORT_229_data = 2'h0;
  assign ram_1_MPORT_229_addr = 8'he5;
  assign ram_1_MPORT_229_mask = 1'h1;
  assign ram_1_MPORT_229_en = reset;
  assign ram_1_MPORT_230_data = 2'h0;
  assign ram_1_MPORT_230_addr = 8'he6;
  assign ram_1_MPORT_230_mask = 1'h1;
  assign ram_1_MPORT_230_en = reset;
  assign ram_1_MPORT_231_data = 2'h0;
  assign ram_1_MPORT_231_addr = 8'he7;
  assign ram_1_MPORT_231_mask = 1'h1;
  assign ram_1_MPORT_231_en = reset;
  assign ram_1_MPORT_232_data = 2'h0;
  assign ram_1_MPORT_232_addr = 8'he8;
  assign ram_1_MPORT_232_mask = 1'h1;
  assign ram_1_MPORT_232_en = reset;
  assign ram_1_MPORT_233_data = 2'h0;
  assign ram_1_MPORT_233_addr = 8'he9;
  assign ram_1_MPORT_233_mask = 1'h1;
  assign ram_1_MPORT_233_en = reset;
  assign ram_1_MPORT_234_data = 2'h0;
  assign ram_1_MPORT_234_addr = 8'hea;
  assign ram_1_MPORT_234_mask = 1'h1;
  assign ram_1_MPORT_234_en = reset;
  assign ram_1_MPORT_235_data = 2'h0;
  assign ram_1_MPORT_235_addr = 8'heb;
  assign ram_1_MPORT_235_mask = 1'h1;
  assign ram_1_MPORT_235_en = reset;
  assign ram_1_MPORT_236_data = 2'h0;
  assign ram_1_MPORT_236_addr = 8'hec;
  assign ram_1_MPORT_236_mask = 1'h1;
  assign ram_1_MPORT_236_en = reset;
  assign ram_1_MPORT_237_data = 2'h0;
  assign ram_1_MPORT_237_addr = 8'hed;
  assign ram_1_MPORT_237_mask = 1'h1;
  assign ram_1_MPORT_237_en = reset;
  assign ram_1_MPORT_238_data = 2'h0;
  assign ram_1_MPORT_238_addr = 8'hee;
  assign ram_1_MPORT_238_mask = 1'h1;
  assign ram_1_MPORT_238_en = reset;
  assign ram_1_MPORT_239_data = 2'h0;
  assign ram_1_MPORT_239_addr = 8'hef;
  assign ram_1_MPORT_239_mask = 1'h1;
  assign ram_1_MPORT_239_en = reset;
  assign ram_1_MPORT_240_data = 2'h0;
  assign ram_1_MPORT_240_addr = 8'hf0;
  assign ram_1_MPORT_240_mask = 1'h1;
  assign ram_1_MPORT_240_en = reset;
  assign ram_1_MPORT_241_data = 2'h0;
  assign ram_1_MPORT_241_addr = 8'hf1;
  assign ram_1_MPORT_241_mask = 1'h1;
  assign ram_1_MPORT_241_en = reset;
  assign ram_1_MPORT_242_data = 2'h0;
  assign ram_1_MPORT_242_addr = 8'hf2;
  assign ram_1_MPORT_242_mask = 1'h1;
  assign ram_1_MPORT_242_en = reset;
  assign ram_1_MPORT_243_data = 2'h0;
  assign ram_1_MPORT_243_addr = 8'hf3;
  assign ram_1_MPORT_243_mask = 1'h1;
  assign ram_1_MPORT_243_en = reset;
  assign ram_1_MPORT_244_data = 2'h0;
  assign ram_1_MPORT_244_addr = 8'hf4;
  assign ram_1_MPORT_244_mask = 1'h1;
  assign ram_1_MPORT_244_en = reset;
  assign ram_1_MPORT_245_data = 2'h0;
  assign ram_1_MPORT_245_addr = 8'hf5;
  assign ram_1_MPORT_245_mask = 1'h1;
  assign ram_1_MPORT_245_en = reset;
  assign ram_1_MPORT_246_data = 2'h0;
  assign ram_1_MPORT_246_addr = 8'hf6;
  assign ram_1_MPORT_246_mask = 1'h1;
  assign ram_1_MPORT_246_en = reset;
  assign ram_1_MPORT_247_data = 2'h0;
  assign ram_1_MPORT_247_addr = 8'hf7;
  assign ram_1_MPORT_247_mask = 1'h1;
  assign ram_1_MPORT_247_en = reset;
  assign ram_1_MPORT_248_data = 2'h0;
  assign ram_1_MPORT_248_addr = 8'hf8;
  assign ram_1_MPORT_248_mask = 1'h1;
  assign ram_1_MPORT_248_en = reset;
  assign ram_1_MPORT_249_data = 2'h0;
  assign ram_1_MPORT_249_addr = 8'hf9;
  assign ram_1_MPORT_249_mask = 1'h1;
  assign ram_1_MPORT_249_en = reset;
  assign ram_1_MPORT_250_data = 2'h0;
  assign ram_1_MPORT_250_addr = 8'hfa;
  assign ram_1_MPORT_250_mask = 1'h1;
  assign ram_1_MPORT_250_en = reset;
  assign ram_1_MPORT_251_data = 2'h0;
  assign ram_1_MPORT_251_addr = 8'hfb;
  assign ram_1_MPORT_251_mask = 1'h1;
  assign ram_1_MPORT_251_en = reset;
  assign ram_1_MPORT_252_data = 2'h0;
  assign ram_1_MPORT_252_addr = 8'hfc;
  assign ram_1_MPORT_252_mask = 1'h1;
  assign ram_1_MPORT_252_en = reset;
  assign ram_1_MPORT_253_data = 2'h0;
  assign ram_1_MPORT_253_addr = 8'hfd;
  assign ram_1_MPORT_253_mask = 1'h1;
  assign ram_1_MPORT_253_en = reset;
  assign ram_1_MPORT_254_data = 2'h0;
  assign ram_1_MPORT_254_addr = 8'hfe;
  assign ram_1_MPORT_254_mask = 1'h1;
  assign ram_1_MPORT_254_en = reset;
  assign ram_1_MPORT_255_data = 2'h0;
  assign ram_1_MPORT_255_addr = 8'hff;
  assign ram_1_MPORT_255_mask = 1'h1;
  assign ram_1_MPORT_255_en = reset;
  assign ram_1_MPORT_256_data = io_wdata[3:2];
  assign ram_1_MPORT_256_addr = io_addr;
  assign ram_1_MPORT_256_mask = io_wmask[1];
  assign ram_1_MPORT_256_en = io_rw;
  assign ram_2_io_rdata_MPORT_en = ram_2_io_rdata_MPORT_en_pipe_0;
  assign ram_2_io_rdata_MPORT_addr = ram_2_io_rdata_MPORT_addr_pipe_0;
  assign ram_2_io_rdata_MPORT_data = ram_2[ram_2_io_rdata_MPORT_addr]; // @[SRAM.scala 36:26]
  assign ram_2_MPORT_data = 2'h0;
  assign ram_2_MPORT_addr = 8'h0;
  assign ram_2_MPORT_mask = 1'h1;
  assign ram_2_MPORT_en = reset;
  assign ram_2_MPORT_1_data = 2'h0;
  assign ram_2_MPORT_1_addr = 8'h1;
  assign ram_2_MPORT_1_mask = 1'h1;
  assign ram_2_MPORT_1_en = reset;
  assign ram_2_MPORT_2_data = 2'h0;
  assign ram_2_MPORT_2_addr = 8'h2;
  assign ram_2_MPORT_2_mask = 1'h1;
  assign ram_2_MPORT_2_en = reset;
  assign ram_2_MPORT_3_data = 2'h0;
  assign ram_2_MPORT_3_addr = 8'h3;
  assign ram_2_MPORT_3_mask = 1'h1;
  assign ram_2_MPORT_3_en = reset;
  assign ram_2_MPORT_4_data = 2'h0;
  assign ram_2_MPORT_4_addr = 8'h4;
  assign ram_2_MPORT_4_mask = 1'h1;
  assign ram_2_MPORT_4_en = reset;
  assign ram_2_MPORT_5_data = 2'h0;
  assign ram_2_MPORT_5_addr = 8'h5;
  assign ram_2_MPORT_5_mask = 1'h1;
  assign ram_2_MPORT_5_en = reset;
  assign ram_2_MPORT_6_data = 2'h0;
  assign ram_2_MPORT_6_addr = 8'h6;
  assign ram_2_MPORT_6_mask = 1'h1;
  assign ram_2_MPORT_6_en = reset;
  assign ram_2_MPORT_7_data = 2'h0;
  assign ram_2_MPORT_7_addr = 8'h7;
  assign ram_2_MPORT_7_mask = 1'h1;
  assign ram_2_MPORT_7_en = reset;
  assign ram_2_MPORT_8_data = 2'h0;
  assign ram_2_MPORT_8_addr = 8'h8;
  assign ram_2_MPORT_8_mask = 1'h1;
  assign ram_2_MPORT_8_en = reset;
  assign ram_2_MPORT_9_data = 2'h0;
  assign ram_2_MPORT_9_addr = 8'h9;
  assign ram_2_MPORT_9_mask = 1'h1;
  assign ram_2_MPORT_9_en = reset;
  assign ram_2_MPORT_10_data = 2'h0;
  assign ram_2_MPORT_10_addr = 8'ha;
  assign ram_2_MPORT_10_mask = 1'h1;
  assign ram_2_MPORT_10_en = reset;
  assign ram_2_MPORT_11_data = 2'h0;
  assign ram_2_MPORT_11_addr = 8'hb;
  assign ram_2_MPORT_11_mask = 1'h1;
  assign ram_2_MPORT_11_en = reset;
  assign ram_2_MPORT_12_data = 2'h0;
  assign ram_2_MPORT_12_addr = 8'hc;
  assign ram_2_MPORT_12_mask = 1'h1;
  assign ram_2_MPORT_12_en = reset;
  assign ram_2_MPORT_13_data = 2'h0;
  assign ram_2_MPORT_13_addr = 8'hd;
  assign ram_2_MPORT_13_mask = 1'h1;
  assign ram_2_MPORT_13_en = reset;
  assign ram_2_MPORT_14_data = 2'h0;
  assign ram_2_MPORT_14_addr = 8'he;
  assign ram_2_MPORT_14_mask = 1'h1;
  assign ram_2_MPORT_14_en = reset;
  assign ram_2_MPORT_15_data = 2'h0;
  assign ram_2_MPORT_15_addr = 8'hf;
  assign ram_2_MPORT_15_mask = 1'h1;
  assign ram_2_MPORT_15_en = reset;
  assign ram_2_MPORT_16_data = 2'h0;
  assign ram_2_MPORT_16_addr = 8'h10;
  assign ram_2_MPORT_16_mask = 1'h1;
  assign ram_2_MPORT_16_en = reset;
  assign ram_2_MPORT_17_data = 2'h0;
  assign ram_2_MPORT_17_addr = 8'h11;
  assign ram_2_MPORT_17_mask = 1'h1;
  assign ram_2_MPORT_17_en = reset;
  assign ram_2_MPORT_18_data = 2'h0;
  assign ram_2_MPORT_18_addr = 8'h12;
  assign ram_2_MPORT_18_mask = 1'h1;
  assign ram_2_MPORT_18_en = reset;
  assign ram_2_MPORT_19_data = 2'h0;
  assign ram_2_MPORT_19_addr = 8'h13;
  assign ram_2_MPORT_19_mask = 1'h1;
  assign ram_2_MPORT_19_en = reset;
  assign ram_2_MPORT_20_data = 2'h0;
  assign ram_2_MPORT_20_addr = 8'h14;
  assign ram_2_MPORT_20_mask = 1'h1;
  assign ram_2_MPORT_20_en = reset;
  assign ram_2_MPORT_21_data = 2'h0;
  assign ram_2_MPORT_21_addr = 8'h15;
  assign ram_2_MPORT_21_mask = 1'h1;
  assign ram_2_MPORT_21_en = reset;
  assign ram_2_MPORT_22_data = 2'h0;
  assign ram_2_MPORT_22_addr = 8'h16;
  assign ram_2_MPORT_22_mask = 1'h1;
  assign ram_2_MPORT_22_en = reset;
  assign ram_2_MPORT_23_data = 2'h0;
  assign ram_2_MPORT_23_addr = 8'h17;
  assign ram_2_MPORT_23_mask = 1'h1;
  assign ram_2_MPORT_23_en = reset;
  assign ram_2_MPORT_24_data = 2'h0;
  assign ram_2_MPORT_24_addr = 8'h18;
  assign ram_2_MPORT_24_mask = 1'h1;
  assign ram_2_MPORT_24_en = reset;
  assign ram_2_MPORT_25_data = 2'h0;
  assign ram_2_MPORT_25_addr = 8'h19;
  assign ram_2_MPORT_25_mask = 1'h1;
  assign ram_2_MPORT_25_en = reset;
  assign ram_2_MPORT_26_data = 2'h0;
  assign ram_2_MPORT_26_addr = 8'h1a;
  assign ram_2_MPORT_26_mask = 1'h1;
  assign ram_2_MPORT_26_en = reset;
  assign ram_2_MPORT_27_data = 2'h0;
  assign ram_2_MPORT_27_addr = 8'h1b;
  assign ram_2_MPORT_27_mask = 1'h1;
  assign ram_2_MPORT_27_en = reset;
  assign ram_2_MPORT_28_data = 2'h0;
  assign ram_2_MPORT_28_addr = 8'h1c;
  assign ram_2_MPORT_28_mask = 1'h1;
  assign ram_2_MPORT_28_en = reset;
  assign ram_2_MPORT_29_data = 2'h0;
  assign ram_2_MPORT_29_addr = 8'h1d;
  assign ram_2_MPORT_29_mask = 1'h1;
  assign ram_2_MPORT_29_en = reset;
  assign ram_2_MPORT_30_data = 2'h0;
  assign ram_2_MPORT_30_addr = 8'h1e;
  assign ram_2_MPORT_30_mask = 1'h1;
  assign ram_2_MPORT_30_en = reset;
  assign ram_2_MPORT_31_data = 2'h0;
  assign ram_2_MPORT_31_addr = 8'h1f;
  assign ram_2_MPORT_31_mask = 1'h1;
  assign ram_2_MPORT_31_en = reset;
  assign ram_2_MPORT_32_data = 2'h0;
  assign ram_2_MPORT_32_addr = 8'h20;
  assign ram_2_MPORT_32_mask = 1'h1;
  assign ram_2_MPORT_32_en = reset;
  assign ram_2_MPORT_33_data = 2'h0;
  assign ram_2_MPORT_33_addr = 8'h21;
  assign ram_2_MPORT_33_mask = 1'h1;
  assign ram_2_MPORT_33_en = reset;
  assign ram_2_MPORT_34_data = 2'h0;
  assign ram_2_MPORT_34_addr = 8'h22;
  assign ram_2_MPORT_34_mask = 1'h1;
  assign ram_2_MPORT_34_en = reset;
  assign ram_2_MPORT_35_data = 2'h0;
  assign ram_2_MPORT_35_addr = 8'h23;
  assign ram_2_MPORT_35_mask = 1'h1;
  assign ram_2_MPORT_35_en = reset;
  assign ram_2_MPORT_36_data = 2'h0;
  assign ram_2_MPORT_36_addr = 8'h24;
  assign ram_2_MPORT_36_mask = 1'h1;
  assign ram_2_MPORT_36_en = reset;
  assign ram_2_MPORT_37_data = 2'h0;
  assign ram_2_MPORT_37_addr = 8'h25;
  assign ram_2_MPORT_37_mask = 1'h1;
  assign ram_2_MPORT_37_en = reset;
  assign ram_2_MPORT_38_data = 2'h0;
  assign ram_2_MPORT_38_addr = 8'h26;
  assign ram_2_MPORT_38_mask = 1'h1;
  assign ram_2_MPORT_38_en = reset;
  assign ram_2_MPORT_39_data = 2'h0;
  assign ram_2_MPORT_39_addr = 8'h27;
  assign ram_2_MPORT_39_mask = 1'h1;
  assign ram_2_MPORT_39_en = reset;
  assign ram_2_MPORT_40_data = 2'h0;
  assign ram_2_MPORT_40_addr = 8'h28;
  assign ram_2_MPORT_40_mask = 1'h1;
  assign ram_2_MPORT_40_en = reset;
  assign ram_2_MPORT_41_data = 2'h0;
  assign ram_2_MPORT_41_addr = 8'h29;
  assign ram_2_MPORT_41_mask = 1'h1;
  assign ram_2_MPORT_41_en = reset;
  assign ram_2_MPORT_42_data = 2'h0;
  assign ram_2_MPORT_42_addr = 8'h2a;
  assign ram_2_MPORT_42_mask = 1'h1;
  assign ram_2_MPORT_42_en = reset;
  assign ram_2_MPORT_43_data = 2'h0;
  assign ram_2_MPORT_43_addr = 8'h2b;
  assign ram_2_MPORT_43_mask = 1'h1;
  assign ram_2_MPORT_43_en = reset;
  assign ram_2_MPORT_44_data = 2'h0;
  assign ram_2_MPORT_44_addr = 8'h2c;
  assign ram_2_MPORT_44_mask = 1'h1;
  assign ram_2_MPORT_44_en = reset;
  assign ram_2_MPORT_45_data = 2'h0;
  assign ram_2_MPORT_45_addr = 8'h2d;
  assign ram_2_MPORT_45_mask = 1'h1;
  assign ram_2_MPORT_45_en = reset;
  assign ram_2_MPORT_46_data = 2'h0;
  assign ram_2_MPORT_46_addr = 8'h2e;
  assign ram_2_MPORT_46_mask = 1'h1;
  assign ram_2_MPORT_46_en = reset;
  assign ram_2_MPORT_47_data = 2'h0;
  assign ram_2_MPORT_47_addr = 8'h2f;
  assign ram_2_MPORT_47_mask = 1'h1;
  assign ram_2_MPORT_47_en = reset;
  assign ram_2_MPORT_48_data = 2'h0;
  assign ram_2_MPORT_48_addr = 8'h30;
  assign ram_2_MPORT_48_mask = 1'h1;
  assign ram_2_MPORT_48_en = reset;
  assign ram_2_MPORT_49_data = 2'h0;
  assign ram_2_MPORT_49_addr = 8'h31;
  assign ram_2_MPORT_49_mask = 1'h1;
  assign ram_2_MPORT_49_en = reset;
  assign ram_2_MPORT_50_data = 2'h0;
  assign ram_2_MPORT_50_addr = 8'h32;
  assign ram_2_MPORT_50_mask = 1'h1;
  assign ram_2_MPORT_50_en = reset;
  assign ram_2_MPORT_51_data = 2'h0;
  assign ram_2_MPORT_51_addr = 8'h33;
  assign ram_2_MPORT_51_mask = 1'h1;
  assign ram_2_MPORT_51_en = reset;
  assign ram_2_MPORT_52_data = 2'h0;
  assign ram_2_MPORT_52_addr = 8'h34;
  assign ram_2_MPORT_52_mask = 1'h1;
  assign ram_2_MPORT_52_en = reset;
  assign ram_2_MPORT_53_data = 2'h0;
  assign ram_2_MPORT_53_addr = 8'h35;
  assign ram_2_MPORT_53_mask = 1'h1;
  assign ram_2_MPORT_53_en = reset;
  assign ram_2_MPORT_54_data = 2'h0;
  assign ram_2_MPORT_54_addr = 8'h36;
  assign ram_2_MPORT_54_mask = 1'h1;
  assign ram_2_MPORT_54_en = reset;
  assign ram_2_MPORT_55_data = 2'h0;
  assign ram_2_MPORT_55_addr = 8'h37;
  assign ram_2_MPORT_55_mask = 1'h1;
  assign ram_2_MPORT_55_en = reset;
  assign ram_2_MPORT_56_data = 2'h0;
  assign ram_2_MPORT_56_addr = 8'h38;
  assign ram_2_MPORT_56_mask = 1'h1;
  assign ram_2_MPORT_56_en = reset;
  assign ram_2_MPORT_57_data = 2'h0;
  assign ram_2_MPORT_57_addr = 8'h39;
  assign ram_2_MPORT_57_mask = 1'h1;
  assign ram_2_MPORT_57_en = reset;
  assign ram_2_MPORT_58_data = 2'h0;
  assign ram_2_MPORT_58_addr = 8'h3a;
  assign ram_2_MPORT_58_mask = 1'h1;
  assign ram_2_MPORT_58_en = reset;
  assign ram_2_MPORT_59_data = 2'h0;
  assign ram_2_MPORT_59_addr = 8'h3b;
  assign ram_2_MPORT_59_mask = 1'h1;
  assign ram_2_MPORT_59_en = reset;
  assign ram_2_MPORT_60_data = 2'h0;
  assign ram_2_MPORT_60_addr = 8'h3c;
  assign ram_2_MPORT_60_mask = 1'h1;
  assign ram_2_MPORT_60_en = reset;
  assign ram_2_MPORT_61_data = 2'h0;
  assign ram_2_MPORT_61_addr = 8'h3d;
  assign ram_2_MPORT_61_mask = 1'h1;
  assign ram_2_MPORT_61_en = reset;
  assign ram_2_MPORT_62_data = 2'h0;
  assign ram_2_MPORT_62_addr = 8'h3e;
  assign ram_2_MPORT_62_mask = 1'h1;
  assign ram_2_MPORT_62_en = reset;
  assign ram_2_MPORT_63_data = 2'h0;
  assign ram_2_MPORT_63_addr = 8'h3f;
  assign ram_2_MPORT_63_mask = 1'h1;
  assign ram_2_MPORT_63_en = reset;
  assign ram_2_MPORT_64_data = 2'h0;
  assign ram_2_MPORT_64_addr = 8'h40;
  assign ram_2_MPORT_64_mask = 1'h1;
  assign ram_2_MPORT_64_en = reset;
  assign ram_2_MPORT_65_data = 2'h0;
  assign ram_2_MPORT_65_addr = 8'h41;
  assign ram_2_MPORT_65_mask = 1'h1;
  assign ram_2_MPORT_65_en = reset;
  assign ram_2_MPORT_66_data = 2'h0;
  assign ram_2_MPORT_66_addr = 8'h42;
  assign ram_2_MPORT_66_mask = 1'h1;
  assign ram_2_MPORT_66_en = reset;
  assign ram_2_MPORT_67_data = 2'h0;
  assign ram_2_MPORT_67_addr = 8'h43;
  assign ram_2_MPORT_67_mask = 1'h1;
  assign ram_2_MPORT_67_en = reset;
  assign ram_2_MPORT_68_data = 2'h0;
  assign ram_2_MPORT_68_addr = 8'h44;
  assign ram_2_MPORT_68_mask = 1'h1;
  assign ram_2_MPORT_68_en = reset;
  assign ram_2_MPORT_69_data = 2'h0;
  assign ram_2_MPORT_69_addr = 8'h45;
  assign ram_2_MPORT_69_mask = 1'h1;
  assign ram_2_MPORT_69_en = reset;
  assign ram_2_MPORT_70_data = 2'h0;
  assign ram_2_MPORT_70_addr = 8'h46;
  assign ram_2_MPORT_70_mask = 1'h1;
  assign ram_2_MPORT_70_en = reset;
  assign ram_2_MPORT_71_data = 2'h0;
  assign ram_2_MPORT_71_addr = 8'h47;
  assign ram_2_MPORT_71_mask = 1'h1;
  assign ram_2_MPORT_71_en = reset;
  assign ram_2_MPORT_72_data = 2'h0;
  assign ram_2_MPORT_72_addr = 8'h48;
  assign ram_2_MPORT_72_mask = 1'h1;
  assign ram_2_MPORT_72_en = reset;
  assign ram_2_MPORT_73_data = 2'h0;
  assign ram_2_MPORT_73_addr = 8'h49;
  assign ram_2_MPORT_73_mask = 1'h1;
  assign ram_2_MPORT_73_en = reset;
  assign ram_2_MPORT_74_data = 2'h0;
  assign ram_2_MPORT_74_addr = 8'h4a;
  assign ram_2_MPORT_74_mask = 1'h1;
  assign ram_2_MPORT_74_en = reset;
  assign ram_2_MPORT_75_data = 2'h0;
  assign ram_2_MPORT_75_addr = 8'h4b;
  assign ram_2_MPORT_75_mask = 1'h1;
  assign ram_2_MPORT_75_en = reset;
  assign ram_2_MPORT_76_data = 2'h0;
  assign ram_2_MPORT_76_addr = 8'h4c;
  assign ram_2_MPORT_76_mask = 1'h1;
  assign ram_2_MPORT_76_en = reset;
  assign ram_2_MPORT_77_data = 2'h0;
  assign ram_2_MPORT_77_addr = 8'h4d;
  assign ram_2_MPORT_77_mask = 1'h1;
  assign ram_2_MPORT_77_en = reset;
  assign ram_2_MPORT_78_data = 2'h0;
  assign ram_2_MPORT_78_addr = 8'h4e;
  assign ram_2_MPORT_78_mask = 1'h1;
  assign ram_2_MPORT_78_en = reset;
  assign ram_2_MPORT_79_data = 2'h0;
  assign ram_2_MPORT_79_addr = 8'h4f;
  assign ram_2_MPORT_79_mask = 1'h1;
  assign ram_2_MPORT_79_en = reset;
  assign ram_2_MPORT_80_data = 2'h0;
  assign ram_2_MPORT_80_addr = 8'h50;
  assign ram_2_MPORT_80_mask = 1'h1;
  assign ram_2_MPORT_80_en = reset;
  assign ram_2_MPORT_81_data = 2'h0;
  assign ram_2_MPORT_81_addr = 8'h51;
  assign ram_2_MPORT_81_mask = 1'h1;
  assign ram_2_MPORT_81_en = reset;
  assign ram_2_MPORT_82_data = 2'h0;
  assign ram_2_MPORT_82_addr = 8'h52;
  assign ram_2_MPORT_82_mask = 1'h1;
  assign ram_2_MPORT_82_en = reset;
  assign ram_2_MPORT_83_data = 2'h0;
  assign ram_2_MPORT_83_addr = 8'h53;
  assign ram_2_MPORT_83_mask = 1'h1;
  assign ram_2_MPORT_83_en = reset;
  assign ram_2_MPORT_84_data = 2'h0;
  assign ram_2_MPORT_84_addr = 8'h54;
  assign ram_2_MPORT_84_mask = 1'h1;
  assign ram_2_MPORT_84_en = reset;
  assign ram_2_MPORT_85_data = 2'h0;
  assign ram_2_MPORT_85_addr = 8'h55;
  assign ram_2_MPORT_85_mask = 1'h1;
  assign ram_2_MPORT_85_en = reset;
  assign ram_2_MPORT_86_data = 2'h0;
  assign ram_2_MPORT_86_addr = 8'h56;
  assign ram_2_MPORT_86_mask = 1'h1;
  assign ram_2_MPORT_86_en = reset;
  assign ram_2_MPORT_87_data = 2'h0;
  assign ram_2_MPORT_87_addr = 8'h57;
  assign ram_2_MPORT_87_mask = 1'h1;
  assign ram_2_MPORT_87_en = reset;
  assign ram_2_MPORT_88_data = 2'h0;
  assign ram_2_MPORT_88_addr = 8'h58;
  assign ram_2_MPORT_88_mask = 1'h1;
  assign ram_2_MPORT_88_en = reset;
  assign ram_2_MPORT_89_data = 2'h0;
  assign ram_2_MPORT_89_addr = 8'h59;
  assign ram_2_MPORT_89_mask = 1'h1;
  assign ram_2_MPORT_89_en = reset;
  assign ram_2_MPORT_90_data = 2'h0;
  assign ram_2_MPORT_90_addr = 8'h5a;
  assign ram_2_MPORT_90_mask = 1'h1;
  assign ram_2_MPORT_90_en = reset;
  assign ram_2_MPORT_91_data = 2'h0;
  assign ram_2_MPORT_91_addr = 8'h5b;
  assign ram_2_MPORT_91_mask = 1'h1;
  assign ram_2_MPORT_91_en = reset;
  assign ram_2_MPORT_92_data = 2'h0;
  assign ram_2_MPORT_92_addr = 8'h5c;
  assign ram_2_MPORT_92_mask = 1'h1;
  assign ram_2_MPORT_92_en = reset;
  assign ram_2_MPORT_93_data = 2'h0;
  assign ram_2_MPORT_93_addr = 8'h5d;
  assign ram_2_MPORT_93_mask = 1'h1;
  assign ram_2_MPORT_93_en = reset;
  assign ram_2_MPORT_94_data = 2'h0;
  assign ram_2_MPORT_94_addr = 8'h5e;
  assign ram_2_MPORT_94_mask = 1'h1;
  assign ram_2_MPORT_94_en = reset;
  assign ram_2_MPORT_95_data = 2'h0;
  assign ram_2_MPORT_95_addr = 8'h5f;
  assign ram_2_MPORT_95_mask = 1'h1;
  assign ram_2_MPORT_95_en = reset;
  assign ram_2_MPORT_96_data = 2'h0;
  assign ram_2_MPORT_96_addr = 8'h60;
  assign ram_2_MPORT_96_mask = 1'h1;
  assign ram_2_MPORT_96_en = reset;
  assign ram_2_MPORT_97_data = 2'h0;
  assign ram_2_MPORT_97_addr = 8'h61;
  assign ram_2_MPORT_97_mask = 1'h1;
  assign ram_2_MPORT_97_en = reset;
  assign ram_2_MPORT_98_data = 2'h0;
  assign ram_2_MPORT_98_addr = 8'h62;
  assign ram_2_MPORT_98_mask = 1'h1;
  assign ram_2_MPORT_98_en = reset;
  assign ram_2_MPORT_99_data = 2'h0;
  assign ram_2_MPORT_99_addr = 8'h63;
  assign ram_2_MPORT_99_mask = 1'h1;
  assign ram_2_MPORT_99_en = reset;
  assign ram_2_MPORT_100_data = 2'h0;
  assign ram_2_MPORT_100_addr = 8'h64;
  assign ram_2_MPORT_100_mask = 1'h1;
  assign ram_2_MPORT_100_en = reset;
  assign ram_2_MPORT_101_data = 2'h0;
  assign ram_2_MPORT_101_addr = 8'h65;
  assign ram_2_MPORT_101_mask = 1'h1;
  assign ram_2_MPORT_101_en = reset;
  assign ram_2_MPORT_102_data = 2'h0;
  assign ram_2_MPORT_102_addr = 8'h66;
  assign ram_2_MPORT_102_mask = 1'h1;
  assign ram_2_MPORT_102_en = reset;
  assign ram_2_MPORT_103_data = 2'h0;
  assign ram_2_MPORT_103_addr = 8'h67;
  assign ram_2_MPORT_103_mask = 1'h1;
  assign ram_2_MPORT_103_en = reset;
  assign ram_2_MPORT_104_data = 2'h0;
  assign ram_2_MPORT_104_addr = 8'h68;
  assign ram_2_MPORT_104_mask = 1'h1;
  assign ram_2_MPORT_104_en = reset;
  assign ram_2_MPORT_105_data = 2'h0;
  assign ram_2_MPORT_105_addr = 8'h69;
  assign ram_2_MPORT_105_mask = 1'h1;
  assign ram_2_MPORT_105_en = reset;
  assign ram_2_MPORT_106_data = 2'h0;
  assign ram_2_MPORT_106_addr = 8'h6a;
  assign ram_2_MPORT_106_mask = 1'h1;
  assign ram_2_MPORT_106_en = reset;
  assign ram_2_MPORT_107_data = 2'h0;
  assign ram_2_MPORT_107_addr = 8'h6b;
  assign ram_2_MPORT_107_mask = 1'h1;
  assign ram_2_MPORT_107_en = reset;
  assign ram_2_MPORT_108_data = 2'h0;
  assign ram_2_MPORT_108_addr = 8'h6c;
  assign ram_2_MPORT_108_mask = 1'h1;
  assign ram_2_MPORT_108_en = reset;
  assign ram_2_MPORT_109_data = 2'h0;
  assign ram_2_MPORT_109_addr = 8'h6d;
  assign ram_2_MPORT_109_mask = 1'h1;
  assign ram_2_MPORT_109_en = reset;
  assign ram_2_MPORT_110_data = 2'h0;
  assign ram_2_MPORT_110_addr = 8'h6e;
  assign ram_2_MPORT_110_mask = 1'h1;
  assign ram_2_MPORT_110_en = reset;
  assign ram_2_MPORT_111_data = 2'h0;
  assign ram_2_MPORT_111_addr = 8'h6f;
  assign ram_2_MPORT_111_mask = 1'h1;
  assign ram_2_MPORT_111_en = reset;
  assign ram_2_MPORT_112_data = 2'h0;
  assign ram_2_MPORT_112_addr = 8'h70;
  assign ram_2_MPORT_112_mask = 1'h1;
  assign ram_2_MPORT_112_en = reset;
  assign ram_2_MPORT_113_data = 2'h0;
  assign ram_2_MPORT_113_addr = 8'h71;
  assign ram_2_MPORT_113_mask = 1'h1;
  assign ram_2_MPORT_113_en = reset;
  assign ram_2_MPORT_114_data = 2'h0;
  assign ram_2_MPORT_114_addr = 8'h72;
  assign ram_2_MPORT_114_mask = 1'h1;
  assign ram_2_MPORT_114_en = reset;
  assign ram_2_MPORT_115_data = 2'h0;
  assign ram_2_MPORT_115_addr = 8'h73;
  assign ram_2_MPORT_115_mask = 1'h1;
  assign ram_2_MPORT_115_en = reset;
  assign ram_2_MPORT_116_data = 2'h0;
  assign ram_2_MPORT_116_addr = 8'h74;
  assign ram_2_MPORT_116_mask = 1'h1;
  assign ram_2_MPORT_116_en = reset;
  assign ram_2_MPORT_117_data = 2'h0;
  assign ram_2_MPORT_117_addr = 8'h75;
  assign ram_2_MPORT_117_mask = 1'h1;
  assign ram_2_MPORT_117_en = reset;
  assign ram_2_MPORT_118_data = 2'h0;
  assign ram_2_MPORT_118_addr = 8'h76;
  assign ram_2_MPORT_118_mask = 1'h1;
  assign ram_2_MPORT_118_en = reset;
  assign ram_2_MPORT_119_data = 2'h0;
  assign ram_2_MPORT_119_addr = 8'h77;
  assign ram_2_MPORT_119_mask = 1'h1;
  assign ram_2_MPORT_119_en = reset;
  assign ram_2_MPORT_120_data = 2'h0;
  assign ram_2_MPORT_120_addr = 8'h78;
  assign ram_2_MPORT_120_mask = 1'h1;
  assign ram_2_MPORT_120_en = reset;
  assign ram_2_MPORT_121_data = 2'h0;
  assign ram_2_MPORT_121_addr = 8'h79;
  assign ram_2_MPORT_121_mask = 1'h1;
  assign ram_2_MPORT_121_en = reset;
  assign ram_2_MPORT_122_data = 2'h0;
  assign ram_2_MPORT_122_addr = 8'h7a;
  assign ram_2_MPORT_122_mask = 1'h1;
  assign ram_2_MPORT_122_en = reset;
  assign ram_2_MPORT_123_data = 2'h0;
  assign ram_2_MPORT_123_addr = 8'h7b;
  assign ram_2_MPORT_123_mask = 1'h1;
  assign ram_2_MPORT_123_en = reset;
  assign ram_2_MPORT_124_data = 2'h0;
  assign ram_2_MPORT_124_addr = 8'h7c;
  assign ram_2_MPORT_124_mask = 1'h1;
  assign ram_2_MPORT_124_en = reset;
  assign ram_2_MPORT_125_data = 2'h0;
  assign ram_2_MPORT_125_addr = 8'h7d;
  assign ram_2_MPORT_125_mask = 1'h1;
  assign ram_2_MPORT_125_en = reset;
  assign ram_2_MPORT_126_data = 2'h0;
  assign ram_2_MPORT_126_addr = 8'h7e;
  assign ram_2_MPORT_126_mask = 1'h1;
  assign ram_2_MPORT_126_en = reset;
  assign ram_2_MPORT_127_data = 2'h0;
  assign ram_2_MPORT_127_addr = 8'h7f;
  assign ram_2_MPORT_127_mask = 1'h1;
  assign ram_2_MPORT_127_en = reset;
  assign ram_2_MPORT_128_data = 2'h0;
  assign ram_2_MPORT_128_addr = 8'h80;
  assign ram_2_MPORT_128_mask = 1'h1;
  assign ram_2_MPORT_128_en = reset;
  assign ram_2_MPORT_129_data = 2'h0;
  assign ram_2_MPORT_129_addr = 8'h81;
  assign ram_2_MPORT_129_mask = 1'h1;
  assign ram_2_MPORT_129_en = reset;
  assign ram_2_MPORT_130_data = 2'h0;
  assign ram_2_MPORT_130_addr = 8'h82;
  assign ram_2_MPORT_130_mask = 1'h1;
  assign ram_2_MPORT_130_en = reset;
  assign ram_2_MPORT_131_data = 2'h0;
  assign ram_2_MPORT_131_addr = 8'h83;
  assign ram_2_MPORT_131_mask = 1'h1;
  assign ram_2_MPORT_131_en = reset;
  assign ram_2_MPORT_132_data = 2'h0;
  assign ram_2_MPORT_132_addr = 8'h84;
  assign ram_2_MPORT_132_mask = 1'h1;
  assign ram_2_MPORT_132_en = reset;
  assign ram_2_MPORT_133_data = 2'h0;
  assign ram_2_MPORT_133_addr = 8'h85;
  assign ram_2_MPORT_133_mask = 1'h1;
  assign ram_2_MPORT_133_en = reset;
  assign ram_2_MPORT_134_data = 2'h0;
  assign ram_2_MPORT_134_addr = 8'h86;
  assign ram_2_MPORT_134_mask = 1'h1;
  assign ram_2_MPORT_134_en = reset;
  assign ram_2_MPORT_135_data = 2'h0;
  assign ram_2_MPORT_135_addr = 8'h87;
  assign ram_2_MPORT_135_mask = 1'h1;
  assign ram_2_MPORT_135_en = reset;
  assign ram_2_MPORT_136_data = 2'h0;
  assign ram_2_MPORT_136_addr = 8'h88;
  assign ram_2_MPORT_136_mask = 1'h1;
  assign ram_2_MPORT_136_en = reset;
  assign ram_2_MPORT_137_data = 2'h0;
  assign ram_2_MPORT_137_addr = 8'h89;
  assign ram_2_MPORT_137_mask = 1'h1;
  assign ram_2_MPORT_137_en = reset;
  assign ram_2_MPORT_138_data = 2'h0;
  assign ram_2_MPORT_138_addr = 8'h8a;
  assign ram_2_MPORT_138_mask = 1'h1;
  assign ram_2_MPORT_138_en = reset;
  assign ram_2_MPORT_139_data = 2'h0;
  assign ram_2_MPORT_139_addr = 8'h8b;
  assign ram_2_MPORT_139_mask = 1'h1;
  assign ram_2_MPORT_139_en = reset;
  assign ram_2_MPORT_140_data = 2'h0;
  assign ram_2_MPORT_140_addr = 8'h8c;
  assign ram_2_MPORT_140_mask = 1'h1;
  assign ram_2_MPORT_140_en = reset;
  assign ram_2_MPORT_141_data = 2'h0;
  assign ram_2_MPORT_141_addr = 8'h8d;
  assign ram_2_MPORT_141_mask = 1'h1;
  assign ram_2_MPORT_141_en = reset;
  assign ram_2_MPORT_142_data = 2'h0;
  assign ram_2_MPORT_142_addr = 8'h8e;
  assign ram_2_MPORT_142_mask = 1'h1;
  assign ram_2_MPORT_142_en = reset;
  assign ram_2_MPORT_143_data = 2'h0;
  assign ram_2_MPORT_143_addr = 8'h8f;
  assign ram_2_MPORT_143_mask = 1'h1;
  assign ram_2_MPORT_143_en = reset;
  assign ram_2_MPORT_144_data = 2'h0;
  assign ram_2_MPORT_144_addr = 8'h90;
  assign ram_2_MPORT_144_mask = 1'h1;
  assign ram_2_MPORT_144_en = reset;
  assign ram_2_MPORT_145_data = 2'h0;
  assign ram_2_MPORT_145_addr = 8'h91;
  assign ram_2_MPORT_145_mask = 1'h1;
  assign ram_2_MPORT_145_en = reset;
  assign ram_2_MPORT_146_data = 2'h0;
  assign ram_2_MPORT_146_addr = 8'h92;
  assign ram_2_MPORT_146_mask = 1'h1;
  assign ram_2_MPORT_146_en = reset;
  assign ram_2_MPORT_147_data = 2'h0;
  assign ram_2_MPORT_147_addr = 8'h93;
  assign ram_2_MPORT_147_mask = 1'h1;
  assign ram_2_MPORT_147_en = reset;
  assign ram_2_MPORT_148_data = 2'h0;
  assign ram_2_MPORT_148_addr = 8'h94;
  assign ram_2_MPORT_148_mask = 1'h1;
  assign ram_2_MPORT_148_en = reset;
  assign ram_2_MPORT_149_data = 2'h0;
  assign ram_2_MPORT_149_addr = 8'h95;
  assign ram_2_MPORT_149_mask = 1'h1;
  assign ram_2_MPORT_149_en = reset;
  assign ram_2_MPORT_150_data = 2'h0;
  assign ram_2_MPORT_150_addr = 8'h96;
  assign ram_2_MPORT_150_mask = 1'h1;
  assign ram_2_MPORT_150_en = reset;
  assign ram_2_MPORT_151_data = 2'h0;
  assign ram_2_MPORT_151_addr = 8'h97;
  assign ram_2_MPORT_151_mask = 1'h1;
  assign ram_2_MPORT_151_en = reset;
  assign ram_2_MPORT_152_data = 2'h0;
  assign ram_2_MPORT_152_addr = 8'h98;
  assign ram_2_MPORT_152_mask = 1'h1;
  assign ram_2_MPORT_152_en = reset;
  assign ram_2_MPORT_153_data = 2'h0;
  assign ram_2_MPORT_153_addr = 8'h99;
  assign ram_2_MPORT_153_mask = 1'h1;
  assign ram_2_MPORT_153_en = reset;
  assign ram_2_MPORT_154_data = 2'h0;
  assign ram_2_MPORT_154_addr = 8'h9a;
  assign ram_2_MPORT_154_mask = 1'h1;
  assign ram_2_MPORT_154_en = reset;
  assign ram_2_MPORT_155_data = 2'h0;
  assign ram_2_MPORT_155_addr = 8'h9b;
  assign ram_2_MPORT_155_mask = 1'h1;
  assign ram_2_MPORT_155_en = reset;
  assign ram_2_MPORT_156_data = 2'h0;
  assign ram_2_MPORT_156_addr = 8'h9c;
  assign ram_2_MPORT_156_mask = 1'h1;
  assign ram_2_MPORT_156_en = reset;
  assign ram_2_MPORT_157_data = 2'h0;
  assign ram_2_MPORT_157_addr = 8'h9d;
  assign ram_2_MPORT_157_mask = 1'h1;
  assign ram_2_MPORT_157_en = reset;
  assign ram_2_MPORT_158_data = 2'h0;
  assign ram_2_MPORT_158_addr = 8'h9e;
  assign ram_2_MPORT_158_mask = 1'h1;
  assign ram_2_MPORT_158_en = reset;
  assign ram_2_MPORT_159_data = 2'h0;
  assign ram_2_MPORT_159_addr = 8'h9f;
  assign ram_2_MPORT_159_mask = 1'h1;
  assign ram_2_MPORT_159_en = reset;
  assign ram_2_MPORT_160_data = 2'h0;
  assign ram_2_MPORT_160_addr = 8'ha0;
  assign ram_2_MPORT_160_mask = 1'h1;
  assign ram_2_MPORT_160_en = reset;
  assign ram_2_MPORT_161_data = 2'h0;
  assign ram_2_MPORT_161_addr = 8'ha1;
  assign ram_2_MPORT_161_mask = 1'h1;
  assign ram_2_MPORT_161_en = reset;
  assign ram_2_MPORT_162_data = 2'h0;
  assign ram_2_MPORT_162_addr = 8'ha2;
  assign ram_2_MPORT_162_mask = 1'h1;
  assign ram_2_MPORT_162_en = reset;
  assign ram_2_MPORT_163_data = 2'h0;
  assign ram_2_MPORT_163_addr = 8'ha3;
  assign ram_2_MPORT_163_mask = 1'h1;
  assign ram_2_MPORT_163_en = reset;
  assign ram_2_MPORT_164_data = 2'h0;
  assign ram_2_MPORT_164_addr = 8'ha4;
  assign ram_2_MPORT_164_mask = 1'h1;
  assign ram_2_MPORT_164_en = reset;
  assign ram_2_MPORT_165_data = 2'h0;
  assign ram_2_MPORT_165_addr = 8'ha5;
  assign ram_2_MPORT_165_mask = 1'h1;
  assign ram_2_MPORT_165_en = reset;
  assign ram_2_MPORT_166_data = 2'h0;
  assign ram_2_MPORT_166_addr = 8'ha6;
  assign ram_2_MPORT_166_mask = 1'h1;
  assign ram_2_MPORT_166_en = reset;
  assign ram_2_MPORT_167_data = 2'h0;
  assign ram_2_MPORT_167_addr = 8'ha7;
  assign ram_2_MPORT_167_mask = 1'h1;
  assign ram_2_MPORT_167_en = reset;
  assign ram_2_MPORT_168_data = 2'h0;
  assign ram_2_MPORT_168_addr = 8'ha8;
  assign ram_2_MPORT_168_mask = 1'h1;
  assign ram_2_MPORT_168_en = reset;
  assign ram_2_MPORT_169_data = 2'h0;
  assign ram_2_MPORT_169_addr = 8'ha9;
  assign ram_2_MPORT_169_mask = 1'h1;
  assign ram_2_MPORT_169_en = reset;
  assign ram_2_MPORT_170_data = 2'h0;
  assign ram_2_MPORT_170_addr = 8'haa;
  assign ram_2_MPORT_170_mask = 1'h1;
  assign ram_2_MPORT_170_en = reset;
  assign ram_2_MPORT_171_data = 2'h0;
  assign ram_2_MPORT_171_addr = 8'hab;
  assign ram_2_MPORT_171_mask = 1'h1;
  assign ram_2_MPORT_171_en = reset;
  assign ram_2_MPORT_172_data = 2'h0;
  assign ram_2_MPORT_172_addr = 8'hac;
  assign ram_2_MPORT_172_mask = 1'h1;
  assign ram_2_MPORT_172_en = reset;
  assign ram_2_MPORT_173_data = 2'h0;
  assign ram_2_MPORT_173_addr = 8'had;
  assign ram_2_MPORT_173_mask = 1'h1;
  assign ram_2_MPORT_173_en = reset;
  assign ram_2_MPORT_174_data = 2'h0;
  assign ram_2_MPORT_174_addr = 8'hae;
  assign ram_2_MPORT_174_mask = 1'h1;
  assign ram_2_MPORT_174_en = reset;
  assign ram_2_MPORT_175_data = 2'h0;
  assign ram_2_MPORT_175_addr = 8'haf;
  assign ram_2_MPORT_175_mask = 1'h1;
  assign ram_2_MPORT_175_en = reset;
  assign ram_2_MPORT_176_data = 2'h0;
  assign ram_2_MPORT_176_addr = 8'hb0;
  assign ram_2_MPORT_176_mask = 1'h1;
  assign ram_2_MPORT_176_en = reset;
  assign ram_2_MPORT_177_data = 2'h0;
  assign ram_2_MPORT_177_addr = 8'hb1;
  assign ram_2_MPORT_177_mask = 1'h1;
  assign ram_2_MPORT_177_en = reset;
  assign ram_2_MPORT_178_data = 2'h0;
  assign ram_2_MPORT_178_addr = 8'hb2;
  assign ram_2_MPORT_178_mask = 1'h1;
  assign ram_2_MPORT_178_en = reset;
  assign ram_2_MPORT_179_data = 2'h0;
  assign ram_2_MPORT_179_addr = 8'hb3;
  assign ram_2_MPORT_179_mask = 1'h1;
  assign ram_2_MPORT_179_en = reset;
  assign ram_2_MPORT_180_data = 2'h0;
  assign ram_2_MPORT_180_addr = 8'hb4;
  assign ram_2_MPORT_180_mask = 1'h1;
  assign ram_2_MPORT_180_en = reset;
  assign ram_2_MPORT_181_data = 2'h0;
  assign ram_2_MPORT_181_addr = 8'hb5;
  assign ram_2_MPORT_181_mask = 1'h1;
  assign ram_2_MPORT_181_en = reset;
  assign ram_2_MPORT_182_data = 2'h0;
  assign ram_2_MPORT_182_addr = 8'hb6;
  assign ram_2_MPORT_182_mask = 1'h1;
  assign ram_2_MPORT_182_en = reset;
  assign ram_2_MPORT_183_data = 2'h0;
  assign ram_2_MPORT_183_addr = 8'hb7;
  assign ram_2_MPORT_183_mask = 1'h1;
  assign ram_2_MPORT_183_en = reset;
  assign ram_2_MPORT_184_data = 2'h0;
  assign ram_2_MPORT_184_addr = 8'hb8;
  assign ram_2_MPORT_184_mask = 1'h1;
  assign ram_2_MPORT_184_en = reset;
  assign ram_2_MPORT_185_data = 2'h0;
  assign ram_2_MPORT_185_addr = 8'hb9;
  assign ram_2_MPORT_185_mask = 1'h1;
  assign ram_2_MPORT_185_en = reset;
  assign ram_2_MPORT_186_data = 2'h0;
  assign ram_2_MPORT_186_addr = 8'hba;
  assign ram_2_MPORT_186_mask = 1'h1;
  assign ram_2_MPORT_186_en = reset;
  assign ram_2_MPORT_187_data = 2'h0;
  assign ram_2_MPORT_187_addr = 8'hbb;
  assign ram_2_MPORT_187_mask = 1'h1;
  assign ram_2_MPORT_187_en = reset;
  assign ram_2_MPORT_188_data = 2'h0;
  assign ram_2_MPORT_188_addr = 8'hbc;
  assign ram_2_MPORT_188_mask = 1'h1;
  assign ram_2_MPORT_188_en = reset;
  assign ram_2_MPORT_189_data = 2'h0;
  assign ram_2_MPORT_189_addr = 8'hbd;
  assign ram_2_MPORT_189_mask = 1'h1;
  assign ram_2_MPORT_189_en = reset;
  assign ram_2_MPORT_190_data = 2'h0;
  assign ram_2_MPORT_190_addr = 8'hbe;
  assign ram_2_MPORT_190_mask = 1'h1;
  assign ram_2_MPORT_190_en = reset;
  assign ram_2_MPORT_191_data = 2'h0;
  assign ram_2_MPORT_191_addr = 8'hbf;
  assign ram_2_MPORT_191_mask = 1'h1;
  assign ram_2_MPORT_191_en = reset;
  assign ram_2_MPORT_192_data = 2'h0;
  assign ram_2_MPORT_192_addr = 8'hc0;
  assign ram_2_MPORT_192_mask = 1'h1;
  assign ram_2_MPORT_192_en = reset;
  assign ram_2_MPORT_193_data = 2'h0;
  assign ram_2_MPORT_193_addr = 8'hc1;
  assign ram_2_MPORT_193_mask = 1'h1;
  assign ram_2_MPORT_193_en = reset;
  assign ram_2_MPORT_194_data = 2'h0;
  assign ram_2_MPORT_194_addr = 8'hc2;
  assign ram_2_MPORT_194_mask = 1'h1;
  assign ram_2_MPORT_194_en = reset;
  assign ram_2_MPORT_195_data = 2'h0;
  assign ram_2_MPORT_195_addr = 8'hc3;
  assign ram_2_MPORT_195_mask = 1'h1;
  assign ram_2_MPORT_195_en = reset;
  assign ram_2_MPORT_196_data = 2'h0;
  assign ram_2_MPORT_196_addr = 8'hc4;
  assign ram_2_MPORT_196_mask = 1'h1;
  assign ram_2_MPORT_196_en = reset;
  assign ram_2_MPORT_197_data = 2'h0;
  assign ram_2_MPORT_197_addr = 8'hc5;
  assign ram_2_MPORT_197_mask = 1'h1;
  assign ram_2_MPORT_197_en = reset;
  assign ram_2_MPORT_198_data = 2'h0;
  assign ram_2_MPORT_198_addr = 8'hc6;
  assign ram_2_MPORT_198_mask = 1'h1;
  assign ram_2_MPORT_198_en = reset;
  assign ram_2_MPORT_199_data = 2'h0;
  assign ram_2_MPORT_199_addr = 8'hc7;
  assign ram_2_MPORT_199_mask = 1'h1;
  assign ram_2_MPORT_199_en = reset;
  assign ram_2_MPORT_200_data = 2'h0;
  assign ram_2_MPORT_200_addr = 8'hc8;
  assign ram_2_MPORT_200_mask = 1'h1;
  assign ram_2_MPORT_200_en = reset;
  assign ram_2_MPORT_201_data = 2'h0;
  assign ram_2_MPORT_201_addr = 8'hc9;
  assign ram_2_MPORT_201_mask = 1'h1;
  assign ram_2_MPORT_201_en = reset;
  assign ram_2_MPORT_202_data = 2'h0;
  assign ram_2_MPORT_202_addr = 8'hca;
  assign ram_2_MPORT_202_mask = 1'h1;
  assign ram_2_MPORT_202_en = reset;
  assign ram_2_MPORT_203_data = 2'h0;
  assign ram_2_MPORT_203_addr = 8'hcb;
  assign ram_2_MPORT_203_mask = 1'h1;
  assign ram_2_MPORT_203_en = reset;
  assign ram_2_MPORT_204_data = 2'h0;
  assign ram_2_MPORT_204_addr = 8'hcc;
  assign ram_2_MPORT_204_mask = 1'h1;
  assign ram_2_MPORT_204_en = reset;
  assign ram_2_MPORT_205_data = 2'h0;
  assign ram_2_MPORT_205_addr = 8'hcd;
  assign ram_2_MPORT_205_mask = 1'h1;
  assign ram_2_MPORT_205_en = reset;
  assign ram_2_MPORT_206_data = 2'h0;
  assign ram_2_MPORT_206_addr = 8'hce;
  assign ram_2_MPORT_206_mask = 1'h1;
  assign ram_2_MPORT_206_en = reset;
  assign ram_2_MPORT_207_data = 2'h0;
  assign ram_2_MPORT_207_addr = 8'hcf;
  assign ram_2_MPORT_207_mask = 1'h1;
  assign ram_2_MPORT_207_en = reset;
  assign ram_2_MPORT_208_data = 2'h0;
  assign ram_2_MPORT_208_addr = 8'hd0;
  assign ram_2_MPORT_208_mask = 1'h1;
  assign ram_2_MPORT_208_en = reset;
  assign ram_2_MPORT_209_data = 2'h0;
  assign ram_2_MPORT_209_addr = 8'hd1;
  assign ram_2_MPORT_209_mask = 1'h1;
  assign ram_2_MPORT_209_en = reset;
  assign ram_2_MPORT_210_data = 2'h0;
  assign ram_2_MPORT_210_addr = 8'hd2;
  assign ram_2_MPORT_210_mask = 1'h1;
  assign ram_2_MPORT_210_en = reset;
  assign ram_2_MPORT_211_data = 2'h0;
  assign ram_2_MPORT_211_addr = 8'hd3;
  assign ram_2_MPORT_211_mask = 1'h1;
  assign ram_2_MPORT_211_en = reset;
  assign ram_2_MPORT_212_data = 2'h0;
  assign ram_2_MPORT_212_addr = 8'hd4;
  assign ram_2_MPORT_212_mask = 1'h1;
  assign ram_2_MPORT_212_en = reset;
  assign ram_2_MPORT_213_data = 2'h0;
  assign ram_2_MPORT_213_addr = 8'hd5;
  assign ram_2_MPORT_213_mask = 1'h1;
  assign ram_2_MPORT_213_en = reset;
  assign ram_2_MPORT_214_data = 2'h0;
  assign ram_2_MPORT_214_addr = 8'hd6;
  assign ram_2_MPORT_214_mask = 1'h1;
  assign ram_2_MPORT_214_en = reset;
  assign ram_2_MPORT_215_data = 2'h0;
  assign ram_2_MPORT_215_addr = 8'hd7;
  assign ram_2_MPORT_215_mask = 1'h1;
  assign ram_2_MPORT_215_en = reset;
  assign ram_2_MPORT_216_data = 2'h0;
  assign ram_2_MPORT_216_addr = 8'hd8;
  assign ram_2_MPORT_216_mask = 1'h1;
  assign ram_2_MPORT_216_en = reset;
  assign ram_2_MPORT_217_data = 2'h0;
  assign ram_2_MPORT_217_addr = 8'hd9;
  assign ram_2_MPORT_217_mask = 1'h1;
  assign ram_2_MPORT_217_en = reset;
  assign ram_2_MPORT_218_data = 2'h0;
  assign ram_2_MPORT_218_addr = 8'hda;
  assign ram_2_MPORT_218_mask = 1'h1;
  assign ram_2_MPORT_218_en = reset;
  assign ram_2_MPORT_219_data = 2'h0;
  assign ram_2_MPORT_219_addr = 8'hdb;
  assign ram_2_MPORT_219_mask = 1'h1;
  assign ram_2_MPORT_219_en = reset;
  assign ram_2_MPORT_220_data = 2'h0;
  assign ram_2_MPORT_220_addr = 8'hdc;
  assign ram_2_MPORT_220_mask = 1'h1;
  assign ram_2_MPORT_220_en = reset;
  assign ram_2_MPORT_221_data = 2'h0;
  assign ram_2_MPORT_221_addr = 8'hdd;
  assign ram_2_MPORT_221_mask = 1'h1;
  assign ram_2_MPORT_221_en = reset;
  assign ram_2_MPORT_222_data = 2'h0;
  assign ram_2_MPORT_222_addr = 8'hde;
  assign ram_2_MPORT_222_mask = 1'h1;
  assign ram_2_MPORT_222_en = reset;
  assign ram_2_MPORT_223_data = 2'h0;
  assign ram_2_MPORT_223_addr = 8'hdf;
  assign ram_2_MPORT_223_mask = 1'h1;
  assign ram_2_MPORT_223_en = reset;
  assign ram_2_MPORT_224_data = 2'h0;
  assign ram_2_MPORT_224_addr = 8'he0;
  assign ram_2_MPORT_224_mask = 1'h1;
  assign ram_2_MPORT_224_en = reset;
  assign ram_2_MPORT_225_data = 2'h0;
  assign ram_2_MPORT_225_addr = 8'he1;
  assign ram_2_MPORT_225_mask = 1'h1;
  assign ram_2_MPORT_225_en = reset;
  assign ram_2_MPORT_226_data = 2'h0;
  assign ram_2_MPORT_226_addr = 8'he2;
  assign ram_2_MPORT_226_mask = 1'h1;
  assign ram_2_MPORT_226_en = reset;
  assign ram_2_MPORT_227_data = 2'h0;
  assign ram_2_MPORT_227_addr = 8'he3;
  assign ram_2_MPORT_227_mask = 1'h1;
  assign ram_2_MPORT_227_en = reset;
  assign ram_2_MPORT_228_data = 2'h0;
  assign ram_2_MPORT_228_addr = 8'he4;
  assign ram_2_MPORT_228_mask = 1'h1;
  assign ram_2_MPORT_228_en = reset;
  assign ram_2_MPORT_229_data = 2'h0;
  assign ram_2_MPORT_229_addr = 8'he5;
  assign ram_2_MPORT_229_mask = 1'h1;
  assign ram_2_MPORT_229_en = reset;
  assign ram_2_MPORT_230_data = 2'h0;
  assign ram_2_MPORT_230_addr = 8'he6;
  assign ram_2_MPORT_230_mask = 1'h1;
  assign ram_2_MPORT_230_en = reset;
  assign ram_2_MPORT_231_data = 2'h0;
  assign ram_2_MPORT_231_addr = 8'he7;
  assign ram_2_MPORT_231_mask = 1'h1;
  assign ram_2_MPORT_231_en = reset;
  assign ram_2_MPORT_232_data = 2'h0;
  assign ram_2_MPORT_232_addr = 8'he8;
  assign ram_2_MPORT_232_mask = 1'h1;
  assign ram_2_MPORT_232_en = reset;
  assign ram_2_MPORT_233_data = 2'h0;
  assign ram_2_MPORT_233_addr = 8'he9;
  assign ram_2_MPORT_233_mask = 1'h1;
  assign ram_2_MPORT_233_en = reset;
  assign ram_2_MPORT_234_data = 2'h0;
  assign ram_2_MPORT_234_addr = 8'hea;
  assign ram_2_MPORT_234_mask = 1'h1;
  assign ram_2_MPORT_234_en = reset;
  assign ram_2_MPORT_235_data = 2'h0;
  assign ram_2_MPORT_235_addr = 8'heb;
  assign ram_2_MPORT_235_mask = 1'h1;
  assign ram_2_MPORT_235_en = reset;
  assign ram_2_MPORT_236_data = 2'h0;
  assign ram_2_MPORT_236_addr = 8'hec;
  assign ram_2_MPORT_236_mask = 1'h1;
  assign ram_2_MPORT_236_en = reset;
  assign ram_2_MPORT_237_data = 2'h0;
  assign ram_2_MPORT_237_addr = 8'hed;
  assign ram_2_MPORT_237_mask = 1'h1;
  assign ram_2_MPORT_237_en = reset;
  assign ram_2_MPORT_238_data = 2'h0;
  assign ram_2_MPORT_238_addr = 8'hee;
  assign ram_2_MPORT_238_mask = 1'h1;
  assign ram_2_MPORT_238_en = reset;
  assign ram_2_MPORT_239_data = 2'h0;
  assign ram_2_MPORT_239_addr = 8'hef;
  assign ram_2_MPORT_239_mask = 1'h1;
  assign ram_2_MPORT_239_en = reset;
  assign ram_2_MPORT_240_data = 2'h0;
  assign ram_2_MPORT_240_addr = 8'hf0;
  assign ram_2_MPORT_240_mask = 1'h1;
  assign ram_2_MPORT_240_en = reset;
  assign ram_2_MPORT_241_data = 2'h0;
  assign ram_2_MPORT_241_addr = 8'hf1;
  assign ram_2_MPORT_241_mask = 1'h1;
  assign ram_2_MPORT_241_en = reset;
  assign ram_2_MPORT_242_data = 2'h0;
  assign ram_2_MPORT_242_addr = 8'hf2;
  assign ram_2_MPORT_242_mask = 1'h1;
  assign ram_2_MPORT_242_en = reset;
  assign ram_2_MPORT_243_data = 2'h0;
  assign ram_2_MPORT_243_addr = 8'hf3;
  assign ram_2_MPORT_243_mask = 1'h1;
  assign ram_2_MPORT_243_en = reset;
  assign ram_2_MPORT_244_data = 2'h0;
  assign ram_2_MPORT_244_addr = 8'hf4;
  assign ram_2_MPORT_244_mask = 1'h1;
  assign ram_2_MPORT_244_en = reset;
  assign ram_2_MPORT_245_data = 2'h0;
  assign ram_2_MPORT_245_addr = 8'hf5;
  assign ram_2_MPORT_245_mask = 1'h1;
  assign ram_2_MPORT_245_en = reset;
  assign ram_2_MPORT_246_data = 2'h0;
  assign ram_2_MPORT_246_addr = 8'hf6;
  assign ram_2_MPORT_246_mask = 1'h1;
  assign ram_2_MPORT_246_en = reset;
  assign ram_2_MPORT_247_data = 2'h0;
  assign ram_2_MPORT_247_addr = 8'hf7;
  assign ram_2_MPORT_247_mask = 1'h1;
  assign ram_2_MPORT_247_en = reset;
  assign ram_2_MPORT_248_data = 2'h0;
  assign ram_2_MPORT_248_addr = 8'hf8;
  assign ram_2_MPORT_248_mask = 1'h1;
  assign ram_2_MPORT_248_en = reset;
  assign ram_2_MPORT_249_data = 2'h0;
  assign ram_2_MPORT_249_addr = 8'hf9;
  assign ram_2_MPORT_249_mask = 1'h1;
  assign ram_2_MPORT_249_en = reset;
  assign ram_2_MPORT_250_data = 2'h0;
  assign ram_2_MPORT_250_addr = 8'hfa;
  assign ram_2_MPORT_250_mask = 1'h1;
  assign ram_2_MPORT_250_en = reset;
  assign ram_2_MPORT_251_data = 2'h0;
  assign ram_2_MPORT_251_addr = 8'hfb;
  assign ram_2_MPORT_251_mask = 1'h1;
  assign ram_2_MPORT_251_en = reset;
  assign ram_2_MPORT_252_data = 2'h0;
  assign ram_2_MPORT_252_addr = 8'hfc;
  assign ram_2_MPORT_252_mask = 1'h1;
  assign ram_2_MPORT_252_en = reset;
  assign ram_2_MPORT_253_data = 2'h0;
  assign ram_2_MPORT_253_addr = 8'hfd;
  assign ram_2_MPORT_253_mask = 1'h1;
  assign ram_2_MPORT_253_en = reset;
  assign ram_2_MPORT_254_data = 2'h0;
  assign ram_2_MPORT_254_addr = 8'hfe;
  assign ram_2_MPORT_254_mask = 1'h1;
  assign ram_2_MPORT_254_en = reset;
  assign ram_2_MPORT_255_data = 2'h0;
  assign ram_2_MPORT_255_addr = 8'hff;
  assign ram_2_MPORT_255_mask = 1'h1;
  assign ram_2_MPORT_255_en = reset;
  assign ram_2_MPORT_256_data = io_wdata[5:4];
  assign ram_2_MPORT_256_addr = io_addr;
  assign ram_2_MPORT_256_mask = io_wmask[2];
  assign ram_2_MPORT_256_en = io_rw;
  assign ram_3_io_rdata_MPORT_en = ram_3_io_rdata_MPORT_en_pipe_0;
  assign ram_3_io_rdata_MPORT_addr = ram_3_io_rdata_MPORT_addr_pipe_0;
  assign ram_3_io_rdata_MPORT_data = ram_3[ram_3_io_rdata_MPORT_addr]; // @[SRAM.scala 36:26]
  assign ram_3_MPORT_data = 2'h0;
  assign ram_3_MPORT_addr = 8'h0;
  assign ram_3_MPORT_mask = 1'h1;
  assign ram_3_MPORT_en = reset;
  assign ram_3_MPORT_1_data = 2'h0;
  assign ram_3_MPORT_1_addr = 8'h1;
  assign ram_3_MPORT_1_mask = 1'h1;
  assign ram_3_MPORT_1_en = reset;
  assign ram_3_MPORT_2_data = 2'h0;
  assign ram_3_MPORT_2_addr = 8'h2;
  assign ram_3_MPORT_2_mask = 1'h1;
  assign ram_3_MPORT_2_en = reset;
  assign ram_3_MPORT_3_data = 2'h0;
  assign ram_3_MPORT_3_addr = 8'h3;
  assign ram_3_MPORT_3_mask = 1'h1;
  assign ram_3_MPORT_3_en = reset;
  assign ram_3_MPORT_4_data = 2'h0;
  assign ram_3_MPORT_4_addr = 8'h4;
  assign ram_3_MPORT_4_mask = 1'h1;
  assign ram_3_MPORT_4_en = reset;
  assign ram_3_MPORT_5_data = 2'h0;
  assign ram_3_MPORT_5_addr = 8'h5;
  assign ram_3_MPORT_5_mask = 1'h1;
  assign ram_3_MPORT_5_en = reset;
  assign ram_3_MPORT_6_data = 2'h0;
  assign ram_3_MPORT_6_addr = 8'h6;
  assign ram_3_MPORT_6_mask = 1'h1;
  assign ram_3_MPORT_6_en = reset;
  assign ram_3_MPORT_7_data = 2'h0;
  assign ram_3_MPORT_7_addr = 8'h7;
  assign ram_3_MPORT_7_mask = 1'h1;
  assign ram_3_MPORT_7_en = reset;
  assign ram_3_MPORT_8_data = 2'h0;
  assign ram_3_MPORT_8_addr = 8'h8;
  assign ram_3_MPORT_8_mask = 1'h1;
  assign ram_3_MPORT_8_en = reset;
  assign ram_3_MPORT_9_data = 2'h0;
  assign ram_3_MPORT_9_addr = 8'h9;
  assign ram_3_MPORT_9_mask = 1'h1;
  assign ram_3_MPORT_9_en = reset;
  assign ram_3_MPORT_10_data = 2'h0;
  assign ram_3_MPORT_10_addr = 8'ha;
  assign ram_3_MPORT_10_mask = 1'h1;
  assign ram_3_MPORT_10_en = reset;
  assign ram_3_MPORT_11_data = 2'h0;
  assign ram_3_MPORT_11_addr = 8'hb;
  assign ram_3_MPORT_11_mask = 1'h1;
  assign ram_3_MPORT_11_en = reset;
  assign ram_3_MPORT_12_data = 2'h0;
  assign ram_3_MPORT_12_addr = 8'hc;
  assign ram_3_MPORT_12_mask = 1'h1;
  assign ram_3_MPORT_12_en = reset;
  assign ram_3_MPORT_13_data = 2'h0;
  assign ram_3_MPORT_13_addr = 8'hd;
  assign ram_3_MPORT_13_mask = 1'h1;
  assign ram_3_MPORT_13_en = reset;
  assign ram_3_MPORT_14_data = 2'h0;
  assign ram_3_MPORT_14_addr = 8'he;
  assign ram_3_MPORT_14_mask = 1'h1;
  assign ram_3_MPORT_14_en = reset;
  assign ram_3_MPORT_15_data = 2'h0;
  assign ram_3_MPORT_15_addr = 8'hf;
  assign ram_3_MPORT_15_mask = 1'h1;
  assign ram_3_MPORT_15_en = reset;
  assign ram_3_MPORT_16_data = 2'h0;
  assign ram_3_MPORT_16_addr = 8'h10;
  assign ram_3_MPORT_16_mask = 1'h1;
  assign ram_3_MPORT_16_en = reset;
  assign ram_3_MPORT_17_data = 2'h0;
  assign ram_3_MPORT_17_addr = 8'h11;
  assign ram_3_MPORT_17_mask = 1'h1;
  assign ram_3_MPORT_17_en = reset;
  assign ram_3_MPORT_18_data = 2'h0;
  assign ram_3_MPORT_18_addr = 8'h12;
  assign ram_3_MPORT_18_mask = 1'h1;
  assign ram_3_MPORT_18_en = reset;
  assign ram_3_MPORT_19_data = 2'h0;
  assign ram_3_MPORT_19_addr = 8'h13;
  assign ram_3_MPORT_19_mask = 1'h1;
  assign ram_3_MPORT_19_en = reset;
  assign ram_3_MPORT_20_data = 2'h0;
  assign ram_3_MPORT_20_addr = 8'h14;
  assign ram_3_MPORT_20_mask = 1'h1;
  assign ram_3_MPORT_20_en = reset;
  assign ram_3_MPORT_21_data = 2'h0;
  assign ram_3_MPORT_21_addr = 8'h15;
  assign ram_3_MPORT_21_mask = 1'h1;
  assign ram_3_MPORT_21_en = reset;
  assign ram_3_MPORT_22_data = 2'h0;
  assign ram_3_MPORT_22_addr = 8'h16;
  assign ram_3_MPORT_22_mask = 1'h1;
  assign ram_3_MPORT_22_en = reset;
  assign ram_3_MPORT_23_data = 2'h0;
  assign ram_3_MPORT_23_addr = 8'h17;
  assign ram_3_MPORT_23_mask = 1'h1;
  assign ram_3_MPORT_23_en = reset;
  assign ram_3_MPORT_24_data = 2'h0;
  assign ram_3_MPORT_24_addr = 8'h18;
  assign ram_3_MPORT_24_mask = 1'h1;
  assign ram_3_MPORT_24_en = reset;
  assign ram_3_MPORT_25_data = 2'h0;
  assign ram_3_MPORT_25_addr = 8'h19;
  assign ram_3_MPORT_25_mask = 1'h1;
  assign ram_3_MPORT_25_en = reset;
  assign ram_3_MPORT_26_data = 2'h0;
  assign ram_3_MPORT_26_addr = 8'h1a;
  assign ram_3_MPORT_26_mask = 1'h1;
  assign ram_3_MPORT_26_en = reset;
  assign ram_3_MPORT_27_data = 2'h0;
  assign ram_3_MPORT_27_addr = 8'h1b;
  assign ram_3_MPORT_27_mask = 1'h1;
  assign ram_3_MPORT_27_en = reset;
  assign ram_3_MPORT_28_data = 2'h0;
  assign ram_3_MPORT_28_addr = 8'h1c;
  assign ram_3_MPORT_28_mask = 1'h1;
  assign ram_3_MPORT_28_en = reset;
  assign ram_3_MPORT_29_data = 2'h0;
  assign ram_3_MPORT_29_addr = 8'h1d;
  assign ram_3_MPORT_29_mask = 1'h1;
  assign ram_3_MPORT_29_en = reset;
  assign ram_3_MPORT_30_data = 2'h0;
  assign ram_3_MPORT_30_addr = 8'h1e;
  assign ram_3_MPORT_30_mask = 1'h1;
  assign ram_3_MPORT_30_en = reset;
  assign ram_3_MPORT_31_data = 2'h0;
  assign ram_3_MPORT_31_addr = 8'h1f;
  assign ram_3_MPORT_31_mask = 1'h1;
  assign ram_3_MPORT_31_en = reset;
  assign ram_3_MPORT_32_data = 2'h0;
  assign ram_3_MPORT_32_addr = 8'h20;
  assign ram_3_MPORT_32_mask = 1'h1;
  assign ram_3_MPORT_32_en = reset;
  assign ram_3_MPORT_33_data = 2'h0;
  assign ram_3_MPORT_33_addr = 8'h21;
  assign ram_3_MPORT_33_mask = 1'h1;
  assign ram_3_MPORT_33_en = reset;
  assign ram_3_MPORT_34_data = 2'h0;
  assign ram_3_MPORT_34_addr = 8'h22;
  assign ram_3_MPORT_34_mask = 1'h1;
  assign ram_3_MPORT_34_en = reset;
  assign ram_3_MPORT_35_data = 2'h0;
  assign ram_3_MPORT_35_addr = 8'h23;
  assign ram_3_MPORT_35_mask = 1'h1;
  assign ram_3_MPORT_35_en = reset;
  assign ram_3_MPORT_36_data = 2'h0;
  assign ram_3_MPORT_36_addr = 8'h24;
  assign ram_3_MPORT_36_mask = 1'h1;
  assign ram_3_MPORT_36_en = reset;
  assign ram_3_MPORT_37_data = 2'h0;
  assign ram_3_MPORT_37_addr = 8'h25;
  assign ram_3_MPORT_37_mask = 1'h1;
  assign ram_3_MPORT_37_en = reset;
  assign ram_3_MPORT_38_data = 2'h0;
  assign ram_3_MPORT_38_addr = 8'h26;
  assign ram_3_MPORT_38_mask = 1'h1;
  assign ram_3_MPORT_38_en = reset;
  assign ram_3_MPORT_39_data = 2'h0;
  assign ram_3_MPORT_39_addr = 8'h27;
  assign ram_3_MPORT_39_mask = 1'h1;
  assign ram_3_MPORT_39_en = reset;
  assign ram_3_MPORT_40_data = 2'h0;
  assign ram_3_MPORT_40_addr = 8'h28;
  assign ram_3_MPORT_40_mask = 1'h1;
  assign ram_3_MPORT_40_en = reset;
  assign ram_3_MPORT_41_data = 2'h0;
  assign ram_3_MPORT_41_addr = 8'h29;
  assign ram_3_MPORT_41_mask = 1'h1;
  assign ram_3_MPORT_41_en = reset;
  assign ram_3_MPORT_42_data = 2'h0;
  assign ram_3_MPORT_42_addr = 8'h2a;
  assign ram_3_MPORT_42_mask = 1'h1;
  assign ram_3_MPORT_42_en = reset;
  assign ram_3_MPORT_43_data = 2'h0;
  assign ram_3_MPORT_43_addr = 8'h2b;
  assign ram_3_MPORT_43_mask = 1'h1;
  assign ram_3_MPORT_43_en = reset;
  assign ram_3_MPORT_44_data = 2'h0;
  assign ram_3_MPORT_44_addr = 8'h2c;
  assign ram_3_MPORT_44_mask = 1'h1;
  assign ram_3_MPORT_44_en = reset;
  assign ram_3_MPORT_45_data = 2'h0;
  assign ram_3_MPORT_45_addr = 8'h2d;
  assign ram_3_MPORT_45_mask = 1'h1;
  assign ram_3_MPORT_45_en = reset;
  assign ram_3_MPORT_46_data = 2'h0;
  assign ram_3_MPORT_46_addr = 8'h2e;
  assign ram_3_MPORT_46_mask = 1'h1;
  assign ram_3_MPORT_46_en = reset;
  assign ram_3_MPORT_47_data = 2'h0;
  assign ram_3_MPORT_47_addr = 8'h2f;
  assign ram_3_MPORT_47_mask = 1'h1;
  assign ram_3_MPORT_47_en = reset;
  assign ram_3_MPORT_48_data = 2'h0;
  assign ram_3_MPORT_48_addr = 8'h30;
  assign ram_3_MPORT_48_mask = 1'h1;
  assign ram_3_MPORT_48_en = reset;
  assign ram_3_MPORT_49_data = 2'h0;
  assign ram_3_MPORT_49_addr = 8'h31;
  assign ram_3_MPORT_49_mask = 1'h1;
  assign ram_3_MPORT_49_en = reset;
  assign ram_3_MPORT_50_data = 2'h0;
  assign ram_3_MPORT_50_addr = 8'h32;
  assign ram_3_MPORT_50_mask = 1'h1;
  assign ram_3_MPORT_50_en = reset;
  assign ram_3_MPORT_51_data = 2'h0;
  assign ram_3_MPORT_51_addr = 8'h33;
  assign ram_3_MPORT_51_mask = 1'h1;
  assign ram_3_MPORT_51_en = reset;
  assign ram_3_MPORT_52_data = 2'h0;
  assign ram_3_MPORT_52_addr = 8'h34;
  assign ram_3_MPORT_52_mask = 1'h1;
  assign ram_3_MPORT_52_en = reset;
  assign ram_3_MPORT_53_data = 2'h0;
  assign ram_3_MPORT_53_addr = 8'h35;
  assign ram_3_MPORT_53_mask = 1'h1;
  assign ram_3_MPORT_53_en = reset;
  assign ram_3_MPORT_54_data = 2'h0;
  assign ram_3_MPORT_54_addr = 8'h36;
  assign ram_3_MPORT_54_mask = 1'h1;
  assign ram_3_MPORT_54_en = reset;
  assign ram_3_MPORT_55_data = 2'h0;
  assign ram_3_MPORT_55_addr = 8'h37;
  assign ram_3_MPORT_55_mask = 1'h1;
  assign ram_3_MPORT_55_en = reset;
  assign ram_3_MPORT_56_data = 2'h0;
  assign ram_3_MPORT_56_addr = 8'h38;
  assign ram_3_MPORT_56_mask = 1'h1;
  assign ram_3_MPORT_56_en = reset;
  assign ram_3_MPORT_57_data = 2'h0;
  assign ram_3_MPORT_57_addr = 8'h39;
  assign ram_3_MPORT_57_mask = 1'h1;
  assign ram_3_MPORT_57_en = reset;
  assign ram_3_MPORT_58_data = 2'h0;
  assign ram_3_MPORT_58_addr = 8'h3a;
  assign ram_3_MPORT_58_mask = 1'h1;
  assign ram_3_MPORT_58_en = reset;
  assign ram_3_MPORT_59_data = 2'h0;
  assign ram_3_MPORT_59_addr = 8'h3b;
  assign ram_3_MPORT_59_mask = 1'h1;
  assign ram_3_MPORT_59_en = reset;
  assign ram_3_MPORT_60_data = 2'h0;
  assign ram_3_MPORT_60_addr = 8'h3c;
  assign ram_3_MPORT_60_mask = 1'h1;
  assign ram_3_MPORT_60_en = reset;
  assign ram_3_MPORT_61_data = 2'h0;
  assign ram_3_MPORT_61_addr = 8'h3d;
  assign ram_3_MPORT_61_mask = 1'h1;
  assign ram_3_MPORT_61_en = reset;
  assign ram_3_MPORT_62_data = 2'h0;
  assign ram_3_MPORT_62_addr = 8'h3e;
  assign ram_3_MPORT_62_mask = 1'h1;
  assign ram_3_MPORT_62_en = reset;
  assign ram_3_MPORT_63_data = 2'h0;
  assign ram_3_MPORT_63_addr = 8'h3f;
  assign ram_3_MPORT_63_mask = 1'h1;
  assign ram_3_MPORT_63_en = reset;
  assign ram_3_MPORT_64_data = 2'h0;
  assign ram_3_MPORT_64_addr = 8'h40;
  assign ram_3_MPORT_64_mask = 1'h1;
  assign ram_3_MPORT_64_en = reset;
  assign ram_3_MPORT_65_data = 2'h0;
  assign ram_3_MPORT_65_addr = 8'h41;
  assign ram_3_MPORT_65_mask = 1'h1;
  assign ram_3_MPORT_65_en = reset;
  assign ram_3_MPORT_66_data = 2'h0;
  assign ram_3_MPORT_66_addr = 8'h42;
  assign ram_3_MPORT_66_mask = 1'h1;
  assign ram_3_MPORT_66_en = reset;
  assign ram_3_MPORT_67_data = 2'h0;
  assign ram_3_MPORT_67_addr = 8'h43;
  assign ram_3_MPORT_67_mask = 1'h1;
  assign ram_3_MPORT_67_en = reset;
  assign ram_3_MPORT_68_data = 2'h0;
  assign ram_3_MPORT_68_addr = 8'h44;
  assign ram_3_MPORT_68_mask = 1'h1;
  assign ram_3_MPORT_68_en = reset;
  assign ram_3_MPORT_69_data = 2'h0;
  assign ram_3_MPORT_69_addr = 8'h45;
  assign ram_3_MPORT_69_mask = 1'h1;
  assign ram_3_MPORT_69_en = reset;
  assign ram_3_MPORT_70_data = 2'h0;
  assign ram_3_MPORT_70_addr = 8'h46;
  assign ram_3_MPORT_70_mask = 1'h1;
  assign ram_3_MPORT_70_en = reset;
  assign ram_3_MPORT_71_data = 2'h0;
  assign ram_3_MPORT_71_addr = 8'h47;
  assign ram_3_MPORT_71_mask = 1'h1;
  assign ram_3_MPORT_71_en = reset;
  assign ram_3_MPORT_72_data = 2'h0;
  assign ram_3_MPORT_72_addr = 8'h48;
  assign ram_3_MPORT_72_mask = 1'h1;
  assign ram_3_MPORT_72_en = reset;
  assign ram_3_MPORT_73_data = 2'h0;
  assign ram_3_MPORT_73_addr = 8'h49;
  assign ram_3_MPORT_73_mask = 1'h1;
  assign ram_3_MPORT_73_en = reset;
  assign ram_3_MPORT_74_data = 2'h0;
  assign ram_3_MPORT_74_addr = 8'h4a;
  assign ram_3_MPORT_74_mask = 1'h1;
  assign ram_3_MPORT_74_en = reset;
  assign ram_3_MPORT_75_data = 2'h0;
  assign ram_3_MPORT_75_addr = 8'h4b;
  assign ram_3_MPORT_75_mask = 1'h1;
  assign ram_3_MPORT_75_en = reset;
  assign ram_3_MPORT_76_data = 2'h0;
  assign ram_3_MPORT_76_addr = 8'h4c;
  assign ram_3_MPORT_76_mask = 1'h1;
  assign ram_3_MPORT_76_en = reset;
  assign ram_3_MPORT_77_data = 2'h0;
  assign ram_3_MPORT_77_addr = 8'h4d;
  assign ram_3_MPORT_77_mask = 1'h1;
  assign ram_3_MPORT_77_en = reset;
  assign ram_3_MPORT_78_data = 2'h0;
  assign ram_3_MPORT_78_addr = 8'h4e;
  assign ram_3_MPORT_78_mask = 1'h1;
  assign ram_3_MPORT_78_en = reset;
  assign ram_3_MPORT_79_data = 2'h0;
  assign ram_3_MPORT_79_addr = 8'h4f;
  assign ram_3_MPORT_79_mask = 1'h1;
  assign ram_3_MPORT_79_en = reset;
  assign ram_3_MPORT_80_data = 2'h0;
  assign ram_3_MPORT_80_addr = 8'h50;
  assign ram_3_MPORT_80_mask = 1'h1;
  assign ram_3_MPORT_80_en = reset;
  assign ram_3_MPORT_81_data = 2'h0;
  assign ram_3_MPORT_81_addr = 8'h51;
  assign ram_3_MPORT_81_mask = 1'h1;
  assign ram_3_MPORT_81_en = reset;
  assign ram_3_MPORT_82_data = 2'h0;
  assign ram_3_MPORT_82_addr = 8'h52;
  assign ram_3_MPORT_82_mask = 1'h1;
  assign ram_3_MPORT_82_en = reset;
  assign ram_3_MPORT_83_data = 2'h0;
  assign ram_3_MPORT_83_addr = 8'h53;
  assign ram_3_MPORT_83_mask = 1'h1;
  assign ram_3_MPORT_83_en = reset;
  assign ram_3_MPORT_84_data = 2'h0;
  assign ram_3_MPORT_84_addr = 8'h54;
  assign ram_3_MPORT_84_mask = 1'h1;
  assign ram_3_MPORT_84_en = reset;
  assign ram_3_MPORT_85_data = 2'h0;
  assign ram_3_MPORT_85_addr = 8'h55;
  assign ram_3_MPORT_85_mask = 1'h1;
  assign ram_3_MPORT_85_en = reset;
  assign ram_3_MPORT_86_data = 2'h0;
  assign ram_3_MPORT_86_addr = 8'h56;
  assign ram_3_MPORT_86_mask = 1'h1;
  assign ram_3_MPORT_86_en = reset;
  assign ram_3_MPORT_87_data = 2'h0;
  assign ram_3_MPORT_87_addr = 8'h57;
  assign ram_3_MPORT_87_mask = 1'h1;
  assign ram_3_MPORT_87_en = reset;
  assign ram_3_MPORT_88_data = 2'h0;
  assign ram_3_MPORT_88_addr = 8'h58;
  assign ram_3_MPORT_88_mask = 1'h1;
  assign ram_3_MPORT_88_en = reset;
  assign ram_3_MPORT_89_data = 2'h0;
  assign ram_3_MPORT_89_addr = 8'h59;
  assign ram_3_MPORT_89_mask = 1'h1;
  assign ram_3_MPORT_89_en = reset;
  assign ram_3_MPORT_90_data = 2'h0;
  assign ram_3_MPORT_90_addr = 8'h5a;
  assign ram_3_MPORT_90_mask = 1'h1;
  assign ram_3_MPORT_90_en = reset;
  assign ram_3_MPORT_91_data = 2'h0;
  assign ram_3_MPORT_91_addr = 8'h5b;
  assign ram_3_MPORT_91_mask = 1'h1;
  assign ram_3_MPORT_91_en = reset;
  assign ram_3_MPORT_92_data = 2'h0;
  assign ram_3_MPORT_92_addr = 8'h5c;
  assign ram_3_MPORT_92_mask = 1'h1;
  assign ram_3_MPORT_92_en = reset;
  assign ram_3_MPORT_93_data = 2'h0;
  assign ram_3_MPORT_93_addr = 8'h5d;
  assign ram_3_MPORT_93_mask = 1'h1;
  assign ram_3_MPORT_93_en = reset;
  assign ram_3_MPORT_94_data = 2'h0;
  assign ram_3_MPORT_94_addr = 8'h5e;
  assign ram_3_MPORT_94_mask = 1'h1;
  assign ram_3_MPORT_94_en = reset;
  assign ram_3_MPORT_95_data = 2'h0;
  assign ram_3_MPORT_95_addr = 8'h5f;
  assign ram_3_MPORT_95_mask = 1'h1;
  assign ram_3_MPORT_95_en = reset;
  assign ram_3_MPORT_96_data = 2'h0;
  assign ram_3_MPORT_96_addr = 8'h60;
  assign ram_3_MPORT_96_mask = 1'h1;
  assign ram_3_MPORT_96_en = reset;
  assign ram_3_MPORT_97_data = 2'h0;
  assign ram_3_MPORT_97_addr = 8'h61;
  assign ram_3_MPORT_97_mask = 1'h1;
  assign ram_3_MPORT_97_en = reset;
  assign ram_3_MPORT_98_data = 2'h0;
  assign ram_3_MPORT_98_addr = 8'h62;
  assign ram_3_MPORT_98_mask = 1'h1;
  assign ram_3_MPORT_98_en = reset;
  assign ram_3_MPORT_99_data = 2'h0;
  assign ram_3_MPORT_99_addr = 8'h63;
  assign ram_3_MPORT_99_mask = 1'h1;
  assign ram_3_MPORT_99_en = reset;
  assign ram_3_MPORT_100_data = 2'h0;
  assign ram_3_MPORT_100_addr = 8'h64;
  assign ram_3_MPORT_100_mask = 1'h1;
  assign ram_3_MPORT_100_en = reset;
  assign ram_3_MPORT_101_data = 2'h0;
  assign ram_3_MPORT_101_addr = 8'h65;
  assign ram_3_MPORT_101_mask = 1'h1;
  assign ram_3_MPORT_101_en = reset;
  assign ram_3_MPORT_102_data = 2'h0;
  assign ram_3_MPORT_102_addr = 8'h66;
  assign ram_3_MPORT_102_mask = 1'h1;
  assign ram_3_MPORT_102_en = reset;
  assign ram_3_MPORT_103_data = 2'h0;
  assign ram_3_MPORT_103_addr = 8'h67;
  assign ram_3_MPORT_103_mask = 1'h1;
  assign ram_3_MPORT_103_en = reset;
  assign ram_3_MPORT_104_data = 2'h0;
  assign ram_3_MPORT_104_addr = 8'h68;
  assign ram_3_MPORT_104_mask = 1'h1;
  assign ram_3_MPORT_104_en = reset;
  assign ram_3_MPORT_105_data = 2'h0;
  assign ram_3_MPORT_105_addr = 8'h69;
  assign ram_3_MPORT_105_mask = 1'h1;
  assign ram_3_MPORT_105_en = reset;
  assign ram_3_MPORT_106_data = 2'h0;
  assign ram_3_MPORT_106_addr = 8'h6a;
  assign ram_3_MPORT_106_mask = 1'h1;
  assign ram_3_MPORT_106_en = reset;
  assign ram_3_MPORT_107_data = 2'h0;
  assign ram_3_MPORT_107_addr = 8'h6b;
  assign ram_3_MPORT_107_mask = 1'h1;
  assign ram_3_MPORT_107_en = reset;
  assign ram_3_MPORT_108_data = 2'h0;
  assign ram_3_MPORT_108_addr = 8'h6c;
  assign ram_3_MPORT_108_mask = 1'h1;
  assign ram_3_MPORT_108_en = reset;
  assign ram_3_MPORT_109_data = 2'h0;
  assign ram_3_MPORT_109_addr = 8'h6d;
  assign ram_3_MPORT_109_mask = 1'h1;
  assign ram_3_MPORT_109_en = reset;
  assign ram_3_MPORT_110_data = 2'h0;
  assign ram_3_MPORT_110_addr = 8'h6e;
  assign ram_3_MPORT_110_mask = 1'h1;
  assign ram_3_MPORT_110_en = reset;
  assign ram_3_MPORT_111_data = 2'h0;
  assign ram_3_MPORT_111_addr = 8'h6f;
  assign ram_3_MPORT_111_mask = 1'h1;
  assign ram_3_MPORT_111_en = reset;
  assign ram_3_MPORT_112_data = 2'h0;
  assign ram_3_MPORT_112_addr = 8'h70;
  assign ram_3_MPORT_112_mask = 1'h1;
  assign ram_3_MPORT_112_en = reset;
  assign ram_3_MPORT_113_data = 2'h0;
  assign ram_3_MPORT_113_addr = 8'h71;
  assign ram_3_MPORT_113_mask = 1'h1;
  assign ram_3_MPORT_113_en = reset;
  assign ram_3_MPORT_114_data = 2'h0;
  assign ram_3_MPORT_114_addr = 8'h72;
  assign ram_3_MPORT_114_mask = 1'h1;
  assign ram_3_MPORT_114_en = reset;
  assign ram_3_MPORT_115_data = 2'h0;
  assign ram_3_MPORT_115_addr = 8'h73;
  assign ram_3_MPORT_115_mask = 1'h1;
  assign ram_3_MPORT_115_en = reset;
  assign ram_3_MPORT_116_data = 2'h0;
  assign ram_3_MPORT_116_addr = 8'h74;
  assign ram_3_MPORT_116_mask = 1'h1;
  assign ram_3_MPORT_116_en = reset;
  assign ram_3_MPORT_117_data = 2'h0;
  assign ram_3_MPORT_117_addr = 8'h75;
  assign ram_3_MPORT_117_mask = 1'h1;
  assign ram_3_MPORT_117_en = reset;
  assign ram_3_MPORT_118_data = 2'h0;
  assign ram_3_MPORT_118_addr = 8'h76;
  assign ram_3_MPORT_118_mask = 1'h1;
  assign ram_3_MPORT_118_en = reset;
  assign ram_3_MPORT_119_data = 2'h0;
  assign ram_3_MPORT_119_addr = 8'h77;
  assign ram_3_MPORT_119_mask = 1'h1;
  assign ram_3_MPORT_119_en = reset;
  assign ram_3_MPORT_120_data = 2'h0;
  assign ram_3_MPORT_120_addr = 8'h78;
  assign ram_3_MPORT_120_mask = 1'h1;
  assign ram_3_MPORT_120_en = reset;
  assign ram_3_MPORT_121_data = 2'h0;
  assign ram_3_MPORT_121_addr = 8'h79;
  assign ram_3_MPORT_121_mask = 1'h1;
  assign ram_3_MPORT_121_en = reset;
  assign ram_3_MPORT_122_data = 2'h0;
  assign ram_3_MPORT_122_addr = 8'h7a;
  assign ram_3_MPORT_122_mask = 1'h1;
  assign ram_3_MPORT_122_en = reset;
  assign ram_3_MPORT_123_data = 2'h0;
  assign ram_3_MPORT_123_addr = 8'h7b;
  assign ram_3_MPORT_123_mask = 1'h1;
  assign ram_3_MPORT_123_en = reset;
  assign ram_3_MPORT_124_data = 2'h0;
  assign ram_3_MPORT_124_addr = 8'h7c;
  assign ram_3_MPORT_124_mask = 1'h1;
  assign ram_3_MPORT_124_en = reset;
  assign ram_3_MPORT_125_data = 2'h0;
  assign ram_3_MPORT_125_addr = 8'h7d;
  assign ram_3_MPORT_125_mask = 1'h1;
  assign ram_3_MPORT_125_en = reset;
  assign ram_3_MPORT_126_data = 2'h0;
  assign ram_3_MPORT_126_addr = 8'h7e;
  assign ram_3_MPORT_126_mask = 1'h1;
  assign ram_3_MPORT_126_en = reset;
  assign ram_3_MPORT_127_data = 2'h0;
  assign ram_3_MPORT_127_addr = 8'h7f;
  assign ram_3_MPORT_127_mask = 1'h1;
  assign ram_3_MPORT_127_en = reset;
  assign ram_3_MPORT_128_data = 2'h0;
  assign ram_3_MPORT_128_addr = 8'h80;
  assign ram_3_MPORT_128_mask = 1'h1;
  assign ram_3_MPORT_128_en = reset;
  assign ram_3_MPORT_129_data = 2'h0;
  assign ram_3_MPORT_129_addr = 8'h81;
  assign ram_3_MPORT_129_mask = 1'h1;
  assign ram_3_MPORT_129_en = reset;
  assign ram_3_MPORT_130_data = 2'h0;
  assign ram_3_MPORT_130_addr = 8'h82;
  assign ram_3_MPORT_130_mask = 1'h1;
  assign ram_3_MPORT_130_en = reset;
  assign ram_3_MPORT_131_data = 2'h0;
  assign ram_3_MPORT_131_addr = 8'h83;
  assign ram_3_MPORT_131_mask = 1'h1;
  assign ram_3_MPORT_131_en = reset;
  assign ram_3_MPORT_132_data = 2'h0;
  assign ram_3_MPORT_132_addr = 8'h84;
  assign ram_3_MPORT_132_mask = 1'h1;
  assign ram_3_MPORT_132_en = reset;
  assign ram_3_MPORT_133_data = 2'h0;
  assign ram_3_MPORT_133_addr = 8'h85;
  assign ram_3_MPORT_133_mask = 1'h1;
  assign ram_3_MPORT_133_en = reset;
  assign ram_3_MPORT_134_data = 2'h0;
  assign ram_3_MPORT_134_addr = 8'h86;
  assign ram_3_MPORT_134_mask = 1'h1;
  assign ram_3_MPORT_134_en = reset;
  assign ram_3_MPORT_135_data = 2'h0;
  assign ram_3_MPORT_135_addr = 8'h87;
  assign ram_3_MPORT_135_mask = 1'h1;
  assign ram_3_MPORT_135_en = reset;
  assign ram_3_MPORT_136_data = 2'h0;
  assign ram_3_MPORT_136_addr = 8'h88;
  assign ram_3_MPORT_136_mask = 1'h1;
  assign ram_3_MPORT_136_en = reset;
  assign ram_3_MPORT_137_data = 2'h0;
  assign ram_3_MPORT_137_addr = 8'h89;
  assign ram_3_MPORT_137_mask = 1'h1;
  assign ram_3_MPORT_137_en = reset;
  assign ram_3_MPORT_138_data = 2'h0;
  assign ram_3_MPORT_138_addr = 8'h8a;
  assign ram_3_MPORT_138_mask = 1'h1;
  assign ram_3_MPORT_138_en = reset;
  assign ram_3_MPORT_139_data = 2'h0;
  assign ram_3_MPORT_139_addr = 8'h8b;
  assign ram_3_MPORT_139_mask = 1'h1;
  assign ram_3_MPORT_139_en = reset;
  assign ram_3_MPORT_140_data = 2'h0;
  assign ram_3_MPORT_140_addr = 8'h8c;
  assign ram_3_MPORT_140_mask = 1'h1;
  assign ram_3_MPORT_140_en = reset;
  assign ram_3_MPORT_141_data = 2'h0;
  assign ram_3_MPORT_141_addr = 8'h8d;
  assign ram_3_MPORT_141_mask = 1'h1;
  assign ram_3_MPORT_141_en = reset;
  assign ram_3_MPORT_142_data = 2'h0;
  assign ram_3_MPORT_142_addr = 8'h8e;
  assign ram_3_MPORT_142_mask = 1'h1;
  assign ram_3_MPORT_142_en = reset;
  assign ram_3_MPORT_143_data = 2'h0;
  assign ram_3_MPORT_143_addr = 8'h8f;
  assign ram_3_MPORT_143_mask = 1'h1;
  assign ram_3_MPORT_143_en = reset;
  assign ram_3_MPORT_144_data = 2'h0;
  assign ram_3_MPORT_144_addr = 8'h90;
  assign ram_3_MPORT_144_mask = 1'h1;
  assign ram_3_MPORT_144_en = reset;
  assign ram_3_MPORT_145_data = 2'h0;
  assign ram_3_MPORT_145_addr = 8'h91;
  assign ram_3_MPORT_145_mask = 1'h1;
  assign ram_3_MPORT_145_en = reset;
  assign ram_3_MPORT_146_data = 2'h0;
  assign ram_3_MPORT_146_addr = 8'h92;
  assign ram_3_MPORT_146_mask = 1'h1;
  assign ram_3_MPORT_146_en = reset;
  assign ram_3_MPORT_147_data = 2'h0;
  assign ram_3_MPORT_147_addr = 8'h93;
  assign ram_3_MPORT_147_mask = 1'h1;
  assign ram_3_MPORT_147_en = reset;
  assign ram_3_MPORT_148_data = 2'h0;
  assign ram_3_MPORT_148_addr = 8'h94;
  assign ram_3_MPORT_148_mask = 1'h1;
  assign ram_3_MPORT_148_en = reset;
  assign ram_3_MPORT_149_data = 2'h0;
  assign ram_3_MPORT_149_addr = 8'h95;
  assign ram_3_MPORT_149_mask = 1'h1;
  assign ram_3_MPORT_149_en = reset;
  assign ram_3_MPORT_150_data = 2'h0;
  assign ram_3_MPORT_150_addr = 8'h96;
  assign ram_3_MPORT_150_mask = 1'h1;
  assign ram_3_MPORT_150_en = reset;
  assign ram_3_MPORT_151_data = 2'h0;
  assign ram_3_MPORT_151_addr = 8'h97;
  assign ram_3_MPORT_151_mask = 1'h1;
  assign ram_3_MPORT_151_en = reset;
  assign ram_3_MPORT_152_data = 2'h0;
  assign ram_3_MPORT_152_addr = 8'h98;
  assign ram_3_MPORT_152_mask = 1'h1;
  assign ram_3_MPORT_152_en = reset;
  assign ram_3_MPORT_153_data = 2'h0;
  assign ram_3_MPORT_153_addr = 8'h99;
  assign ram_3_MPORT_153_mask = 1'h1;
  assign ram_3_MPORT_153_en = reset;
  assign ram_3_MPORT_154_data = 2'h0;
  assign ram_3_MPORT_154_addr = 8'h9a;
  assign ram_3_MPORT_154_mask = 1'h1;
  assign ram_3_MPORT_154_en = reset;
  assign ram_3_MPORT_155_data = 2'h0;
  assign ram_3_MPORT_155_addr = 8'h9b;
  assign ram_3_MPORT_155_mask = 1'h1;
  assign ram_3_MPORT_155_en = reset;
  assign ram_3_MPORT_156_data = 2'h0;
  assign ram_3_MPORT_156_addr = 8'h9c;
  assign ram_3_MPORT_156_mask = 1'h1;
  assign ram_3_MPORT_156_en = reset;
  assign ram_3_MPORT_157_data = 2'h0;
  assign ram_3_MPORT_157_addr = 8'h9d;
  assign ram_3_MPORT_157_mask = 1'h1;
  assign ram_3_MPORT_157_en = reset;
  assign ram_3_MPORT_158_data = 2'h0;
  assign ram_3_MPORT_158_addr = 8'h9e;
  assign ram_3_MPORT_158_mask = 1'h1;
  assign ram_3_MPORT_158_en = reset;
  assign ram_3_MPORT_159_data = 2'h0;
  assign ram_3_MPORT_159_addr = 8'h9f;
  assign ram_3_MPORT_159_mask = 1'h1;
  assign ram_3_MPORT_159_en = reset;
  assign ram_3_MPORT_160_data = 2'h0;
  assign ram_3_MPORT_160_addr = 8'ha0;
  assign ram_3_MPORT_160_mask = 1'h1;
  assign ram_3_MPORT_160_en = reset;
  assign ram_3_MPORT_161_data = 2'h0;
  assign ram_3_MPORT_161_addr = 8'ha1;
  assign ram_3_MPORT_161_mask = 1'h1;
  assign ram_3_MPORT_161_en = reset;
  assign ram_3_MPORT_162_data = 2'h0;
  assign ram_3_MPORT_162_addr = 8'ha2;
  assign ram_3_MPORT_162_mask = 1'h1;
  assign ram_3_MPORT_162_en = reset;
  assign ram_3_MPORT_163_data = 2'h0;
  assign ram_3_MPORT_163_addr = 8'ha3;
  assign ram_3_MPORT_163_mask = 1'h1;
  assign ram_3_MPORT_163_en = reset;
  assign ram_3_MPORT_164_data = 2'h0;
  assign ram_3_MPORT_164_addr = 8'ha4;
  assign ram_3_MPORT_164_mask = 1'h1;
  assign ram_3_MPORT_164_en = reset;
  assign ram_3_MPORT_165_data = 2'h0;
  assign ram_3_MPORT_165_addr = 8'ha5;
  assign ram_3_MPORT_165_mask = 1'h1;
  assign ram_3_MPORT_165_en = reset;
  assign ram_3_MPORT_166_data = 2'h0;
  assign ram_3_MPORT_166_addr = 8'ha6;
  assign ram_3_MPORT_166_mask = 1'h1;
  assign ram_3_MPORT_166_en = reset;
  assign ram_3_MPORT_167_data = 2'h0;
  assign ram_3_MPORT_167_addr = 8'ha7;
  assign ram_3_MPORT_167_mask = 1'h1;
  assign ram_3_MPORT_167_en = reset;
  assign ram_3_MPORT_168_data = 2'h0;
  assign ram_3_MPORT_168_addr = 8'ha8;
  assign ram_3_MPORT_168_mask = 1'h1;
  assign ram_3_MPORT_168_en = reset;
  assign ram_3_MPORT_169_data = 2'h0;
  assign ram_3_MPORT_169_addr = 8'ha9;
  assign ram_3_MPORT_169_mask = 1'h1;
  assign ram_3_MPORT_169_en = reset;
  assign ram_3_MPORT_170_data = 2'h0;
  assign ram_3_MPORT_170_addr = 8'haa;
  assign ram_3_MPORT_170_mask = 1'h1;
  assign ram_3_MPORT_170_en = reset;
  assign ram_3_MPORT_171_data = 2'h0;
  assign ram_3_MPORT_171_addr = 8'hab;
  assign ram_3_MPORT_171_mask = 1'h1;
  assign ram_3_MPORT_171_en = reset;
  assign ram_3_MPORT_172_data = 2'h0;
  assign ram_3_MPORT_172_addr = 8'hac;
  assign ram_3_MPORT_172_mask = 1'h1;
  assign ram_3_MPORT_172_en = reset;
  assign ram_3_MPORT_173_data = 2'h0;
  assign ram_3_MPORT_173_addr = 8'had;
  assign ram_3_MPORT_173_mask = 1'h1;
  assign ram_3_MPORT_173_en = reset;
  assign ram_3_MPORT_174_data = 2'h0;
  assign ram_3_MPORT_174_addr = 8'hae;
  assign ram_3_MPORT_174_mask = 1'h1;
  assign ram_3_MPORT_174_en = reset;
  assign ram_3_MPORT_175_data = 2'h0;
  assign ram_3_MPORT_175_addr = 8'haf;
  assign ram_3_MPORT_175_mask = 1'h1;
  assign ram_3_MPORT_175_en = reset;
  assign ram_3_MPORT_176_data = 2'h0;
  assign ram_3_MPORT_176_addr = 8'hb0;
  assign ram_3_MPORT_176_mask = 1'h1;
  assign ram_3_MPORT_176_en = reset;
  assign ram_3_MPORT_177_data = 2'h0;
  assign ram_3_MPORT_177_addr = 8'hb1;
  assign ram_3_MPORT_177_mask = 1'h1;
  assign ram_3_MPORT_177_en = reset;
  assign ram_3_MPORT_178_data = 2'h0;
  assign ram_3_MPORT_178_addr = 8'hb2;
  assign ram_3_MPORT_178_mask = 1'h1;
  assign ram_3_MPORT_178_en = reset;
  assign ram_3_MPORT_179_data = 2'h0;
  assign ram_3_MPORT_179_addr = 8'hb3;
  assign ram_3_MPORT_179_mask = 1'h1;
  assign ram_3_MPORT_179_en = reset;
  assign ram_3_MPORT_180_data = 2'h0;
  assign ram_3_MPORT_180_addr = 8'hb4;
  assign ram_3_MPORT_180_mask = 1'h1;
  assign ram_3_MPORT_180_en = reset;
  assign ram_3_MPORT_181_data = 2'h0;
  assign ram_3_MPORT_181_addr = 8'hb5;
  assign ram_3_MPORT_181_mask = 1'h1;
  assign ram_3_MPORT_181_en = reset;
  assign ram_3_MPORT_182_data = 2'h0;
  assign ram_3_MPORT_182_addr = 8'hb6;
  assign ram_3_MPORT_182_mask = 1'h1;
  assign ram_3_MPORT_182_en = reset;
  assign ram_3_MPORT_183_data = 2'h0;
  assign ram_3_MPORT_183_addr = 8'hb7;
  assign ram_3_MPORT_183_mask = 1'h1;
  assign ram_3_MPORT_183_en = reset;
  assign ram_3_MPORT_184_data = 2'h0;
  assign ram_3_MPORT_184_addr = 8'hb8;
  assign ram_3_MPORT_184_mask = 1'h1;
  assign ram_3_MPORT_184_en = reset;
  assign ram_3_MPORT_185_data = 2'h0;
  assign ram_3_MPORT_185_addr = 8'hb9;
  assign ram_3_MPORT_185_mask = 1'h1;
  assign ram_3_MPORT_185_en = reset;
  assign ram_3_MPORT_186_data = 2'h0;
  assign ram_3_MPORT_186_addr = 8'hba;
  assign ram_3_MPORT_186_mask = 1'h1;
  assign ram_3_MPORT_186_en = reset;
  assign ram_3_MPORT_187_data = 2'h0;
  assign ram_3_MPORT_187_addr = 8'hbb;
  assign ram_3_MPORT_187_mask = 1'h1;
  assign ram_3_MPORT_187_en = reset;
  assign ram_3_MPORT_188_data = 2'h0;
  assign ram_3_MPORT_188_addr = 8'hbc;
  assign ram_3_MPORT_188_mask = 1'h1;
  assign ram_3_MPORT_188_en = reset;
  assign ram_3_MPORT_189_data = 2'h0;
  assign ram_3_MPORT_189_addr = 8'hbd;
  assign ram_3_MPORT_189_mask = 1'h1;
  assign ram_3_MPORT_189_en = reset;
  assign ram_3_MPORT_190_data = 2'h0;
  assign ram_3_MPORT_190_addr = 8'hbe;
  assign ram_3_MPORT_190_mask = 1'h1;
  assign ram_3_MPORT_190_en = reset;
  assign ram_3_MPORT_191_data = 2'h0;
  assign ram_3_MPORT_191_addr = 8'hbf;
  assign ram_3_MPORT_191_mask = 1'h1;
  assign ram_3_MPORT_191_en = reset;
  assign ram_3_MPORT_192_data = 2'h0;
  assign ram_3_MPORT_192_addr = 8'hc0;
  assign ram_3_MPORT_192_mask = 1'h1;
  assign ram_3_MPORT_192_en = reset;
  assign ram_3_MPORT_193_data = 2'h0;
  assign ram_3_MPORT_193_addr = 8'hc1;
  assign ram_3_MPORT_193_mask = 1'h1;
  assign ram_3_MPORT_193_en = reset;
  assign ram_3_MPORT_194_data = 2'h0;
  assign ram_3_MPORT_194_addr = 8'hc2;
  assign ram_3_MPORT_194_mask = 1'h1;
  assign ram_3_MPORT_194_en = reset;
  assign ram_3_MPORT_195_data = 2'h0;
  assign ram_3_MPORT_195_addr = 8'hc3;
  assign ram_3_MPORT_195_mask = 1'h1;
  assign ram_3_MPORT_195_en = reset;
  assign ram_3_MPORT_196_data = 2'h0;
  assign ram_3_MPORT_196_addr = 8'hc4;
  assign ram_3_MPORT_196_mask = 1'h1;
  assign ram_3_MPORT_196_en = reset;
  assign ram_3_MPORT_197_data = 2'h0;
  assign ram_3_MPORT_197_addr = 8'hc5;
  assign ram_3_MPORT_197_mask = 1'h1;
  assign ram_3_MPORT_197_en = reset;
  assign ram_3_MPORT_198_data = 2'h0;
  assign ram_3_MPORT_198_addr = 8'hc6;
  assign ram_3_MPORT_198_mask = 1'h1;
  assign ram_3_MPORT_198_en = reset;
  assign ram_3_MPORT_199_data = 2'h0;
  assign ram_3_MPORT_199_addr = 8'hc7;
  assign ram_3_MPORT_199_mask = 1'h1;
  assign ram_3_MPORT_199_en = reset;
  assign ram_3_MPORT_200_data = 2'h0;
  assign ram_3_MPORT_200_addr = 8'hc8;
  assign ram_3_MPORT_200_mask = 1'h1;
  assign ram_3_MPORT_200_en = reset;
  assign ram_3_MPORT_201_data = 2'h0;
  assign ram_3_MPORT_201_addr = 8'hc9;
  assign ram_3_MPORT_201_mask = 1'h1;
  assign ram_3_MPORT_201_en = reset;
  assign ram_3_MPORT_202_data = 2'h0;
  assign ram_3_MPORT_202_addr = 8'hca;
  assign ram_3_MPORT_202_mask = 1'h1;
  assign ram_3_MPORT_202_en = reset;
  assign ram_3_MPORT_203_data = 2'h0;
  assign ram_3_MPORT_203_addr = 8'hcb;
  assign ram_3_MPORT_203_mask = 1'h1;
  assign ram_3_MPORT_203_en = reset;
  assign ram_3_MPORT_204_data = 2'h0;
  assign ram_3_MPORT_204_addr = 8'hcc;
  assign ram_3_MPORT_204_mask = 1'h1;
  assign ram_3_MPORT_204_en = reset;
  assign ram_3_MPORT_205_data = 2'h0;
  assign ram_3_MPORT_205_addr = 8'hcd;
  assign ram_3_MPORT_205_mask = 1'h1;
  assign ram_3_MPORT_205_en = reset;
  assign ram_3_MPORT_206_data = 2'h0;
  assign ram_3_MPORT_206_addr = 8'hce;
  assign ram_3_MPORT_206_mask = 1'h1;
  assign ram_3_MPORT_206_en = reset;
  assign ram_3_MPORT_207_data = 2'h0;
  assign ram_3_MPORT_207_addr = 8'hcf;
  assign ram_3_MPORT_207_mask = 1'h1;
  assign ram_3_MPORT_207_en = reset;
  assign ram_3_MPORT_208_data = 2'h0;
  assign ram_3_MPORT_208_addr = 8'hd0;
  assign ram_3_MPORT_208_mask = 1'h1;
  assign ram_3_MPORT_208_en = reset;
  assign ram_3_MPORT_209_data = 2'h0;
  assign ram_3_MPORT_209_addr = 8'hd1;
  assign ram_3_MPORT_209_mask = 1'h1;
  assign ram_3_MPORT_209_en = reset;
  assign ram_3_MPORT_210_data = 2'h0;
  assign ram_3_MPORT_210_addr = 8'hd2;
  assign ram_3_MPORT_210_mask = 1'h1;
  assign ram_3_MPORT_210_en = reset;
  assign ram_3_MPORT_211_data = 2'h0;
  assign ram_3_MPORT_211_addr = 8'hd3;
  assign ram_3_MPORT_211_mask = 1'h1;
  assign ram_3_MPORT_211_en = reset;
  assign ram_3_MPORT_212_data = 2'h0;
  assign ram_3_MPORT_212_addr = 8'hd4;
  assign ram_3_MPORT_212_mask = 1'h1;
  assign ram_3_MPORT_212_en = reset;
  assign ram_3_MPORT_213_data = 2'h0;
  assign ram_3_MPORT_213_addr = 8'hd5;
  assign ram_3_MPORT_213_mask = 1'h1;
  assign ram_3_MPORT_213_en = reset;
  assign ram_3_MPORT_214_data = 2'h0;
  assign ram_3_MPORT_214_addr = 8'hd6;
  assign ram_3_MPORT_214_mask = 1'h1;
  assign ram_3_MPORT_214_en = reset;
  assign ram_3_MPORT_215_data = 2'h0;
  assign ram_3_MPORT_215_addr = 8'hd7;
  assign ram_3_MPORT_215_mask = 1'h1;
  assign ram_3_MPORT_215_en = reset;
  assign ram_3_MPORT_216_data = 2'h0;
  assign ram_3_MPORT_216_addr = 8'hd8;
  assign ram_3_MPORT_216_mask = 1'h1;
  assign ram_3_MPORT_216_en = reset;
  assign ram_3_MPORT_217_data = 2'h0;
  assign ram_3_MPORT_217_addr = 8'hd9;
  assign ram_3_MPORT_217_mask = 1'h1;
  assign ram_3_MPORT_217_en = reset;
  assign ram_3_MPORT_218_data = 2'h0;
  assign ram_3_MPORT_218_addr = 8'hda;
  assign ram_3_MPORT_218_mask = 1'h1;
  assign ram_3_MPORT_218_en = reset;
  assign ram_3_MPORT_219_data = 2'h0;
  assign ram_3_MPORT_219_addr = 8'hdb;
  assign ram_3_MPORT_219_mask = 1'h1;
  assign ram_3_MPORT_219_en = reset;
  assign ram_3_MPORT_220_data = 2'h0;
  assign ram_3_MPORT_220_addr = 8'hdc;
  assign ram_3_MPORT_220_mask = 1'h1;
  assign ram_3_MPORT_220_en = reset;
  assign ram_3_MPORT_221_data = 2'h0;
  assign ram_3_MPORT_221_addr = 8'hdd;
  assign ram_3_MPORT_221_mask = 1'h1;
  assign ram_3_MPORT_221_en = reset;
  assign ram_3_MPORT_222_data = 2'h0;
  assign ram_3_MPORT_222_addr = 8'hde;
  assign ram_3_MPORT_222_mask = 1'h1;
  assign ram_3_MPORT_222_en = reset;
  assign ram_3_MPORT_223_data = 2'h0;
  assign ram_3_MPORT_223_addr = 8'hdf;
  assign ram_3_MPORT_223_mask = 1'h1;
  assign ram_3_MPORT_223_en = reset;
  assign ram_3_MPORT_224_data = 2'h0;
  assign ram_3_MPORT_224_addr = 8'he0;
  assign ram_3_MPORT_224_mask = 1'h1;
  assign ram_3_MPORT_224_en = reset;
  assign ram_3_MPORT_225_data = 2'h0;
  assign ram_3_MPORT_225_addr = 8'he1;
  assign ram_3_MPORT_225_mask = 1'h1;
  assign ram_3_MPORT_225_en = reset;
  assign ram_3_MPORT_226_data = 2'h0;
  assign ram_3_MPORT_226_addr = 8'he2;
  assign ram_3_MPORT_226_mask = 1'h1;
  assign ram_3_MPORT_226_en = reset;
  assign ram_3_MPORT_227_data = 2'h0;
  assign ram_3_MPORT_227_addr = 8'he3;
  assign ram_3_MPORT_227_mask = 1'h1;
  assign ram_3_MPORT_227_en = reset;
  assign ram_3_MPORT_228_data = 2'h0;
  assign ram_3_MPORT_228_addr = 8'he4;
  assign ram_3_MPORT_228_mask = 1'h1;
  assign ram_3_MPORT_228_en = reset;
  assign ram_3_MPORT_229_data = 2'h0;
  assign ram_3_MPORT_229_addr = 8'he5;
  assign ram_3_MPORT_229_mask = 1'h1;
  assign ram_3_MPORT_229_en = reset;
  assign ram_3_MPORT_230_data = 2'h0;
  assign ram_3_MPORT_230_addr = 8'he6;
  assign ram_3_MPORT_230_mask = 1'h1;
  assign ram_3_MPORT_230_en = reset;
  assign ram_3_MPORT_231_data = 2'h0;
  assign ram_3_MPORT_231_addr = 8'he7;
  assign ram_3_MPORT_231_mask = 1'h1;
  assign ram_3_MPORT_231_en = reset;
  assign ram_3_MPORT_232_data = 2'h0;
  assign ram_3_MPORT_232_addr = 8'he8;
  assign ram_3_MPORT_232_mask = 1'h1;
  assign ram_3_MPORT_232_en = reset;
  assign ram_3_MPORT_233_data = 2'h0;
  assign ram_3_MPORT_233_addr = 8'he9;
  assign ram_3_MPORT_233_mask = 1'h1;
  assign ram_3_MPORT_233_en = reset;
  assign ram_3_MPORT_234_data = 2'h0;
  assign ram_3_MPORT_234_addr = 8'hea;
  assign ram_3_MPORT_234_mask = 1'h1;
  assign ram_3_MPORT_234_en = reset;
  assign ram_3_MPORT_235_data = 2'h0;
  assign ram_3_MPORT_235_addr = 8'heb;
  assign ram_3_MPORT_235_mask = 1'h1;
  assign ram_3_MPORT_235_en = reset;
  assign ram_3_MPORT_236_data = 2'h0;
  assign ram_3_MPORT_236_addr = 8'hec;
  assign ram_3_MPORT_236_mask = 1'h1;
  assign ram_3_MPORT_236_en = reset;
  assign ram_3_MPORT_237_data = 2'h0;
  assign ram_3_MPORT_237_addr = 8'hed;
  assign ram_3_MPORT_237_mask = 1'h1;
  assign ram_3_MPORT_237_en = reset;
  assign ram_3_MPORT_238_data = 2'h0;
  assign ram_3_MPORT_238_addr = 8'hee;
  assign ram_3_MPORT_238_mask = 1'h1;
  assign ram_3_MPORT_238_en = reset;
  assign ram_3_MPORT_239_data = 2'h0;
  assign ram_3_MPORT_239_addr = 8'hef;
  assign ram_3_MPORT_239_mask = 1'h1;
  assign ram_3_MPORT_239_en = reset;
  assign ram_3_MPORT_240_data = 2'h0;
  assign ram_3_MPORT_240_addr = 8'hf0;
  assign ram_3_MPORT_240_mask = 1'h1;
  assign ram_3_MPORT_240_en = reset;
  assign ram_3_MPORT_241_data = 2'h0;
  assign ram_3_MPORT_241_addr = 8'hf1;
  assign ram_3_MPORT_241_mask = 1'h1;
  assign ram_3_MPORT_241_en = reset;
  assign ram_3_MPORT_242_data = 2'h0;
  assign ram_3_MPORT_242_addr = 8'hf2;
  assign ram_3_MPORT_242_mask = 1'h1;
  assign ram_3_MPORT_242_en = reset;
  assign ram_3_MPORT_243_data = 2'h0;
  assign ram_3_MPORT_243_addr = 8'hf3;
  assign ram_3_MPORT_243_mask = 1'h1;
  assign ram_3_MPORT_243_en = reset;
  assign ram_3_MPORT_244_data = 2'h0;
  assign ram_3_MPORT_244_addr = 8'hf4;
  assign ram_3_MPORT_244_mask = 1'h1;
  assign ram_3_MPORT_244_en = reset;
  assign ram_3_MPORT_245_data = 2'h0;
  assign ram_3_MPORT_245_addr = 8'hf5;
  assign ram_3_MPORT_245_mask = 1'h1;
  assign ram_3_MPORT_245_en = reset;
  assign ram_3_MPORT_246_data = 2'h0;
  assign ram_3_MPORT_246_addr = 8'hf6;
  assign ram_3_MPORT_246_mask = 1'h1;
  assign ram_3_MPORT_246_en = reset;
  assign ram_3_MPORT_247_data = 2'h0;
  assign ram_3_MPORT_247_addr = 8'hf7;
  assign ram_3_MPORT_247_mask = 1'h1;
  assign ram_3_MPORT_247_en = reset;
  assign ram_3_MPORT_248_data = 2'h0;
  assign ram_3_MPORT_248_addr = 8'hf8;
  assign ram_3_MPORT_248_mask = 1'h1;
  assign ram_3_MPORT_248_en = reset;
  assign ram_3_MPORT_249_data = 2'h0;
  assign ram_3_MPORT_249_addr = 8'hf9;
  assign ram_3_MPORT_249_mask = 1'h1;
  assign ram_3_MPORT_249_en = reset;
  assign ram_3_MPORT_250_data = 2'h0;
  assign ram_3_MPORT_250_addr = 8'hfa;
  assign ram_3_MPORT_250_mask = 1'h1;
  assign ram_3_MPORT_250_en = reset;
  assign ram_3_MPORT_251_data = 2'h0;
  assign ram_3_MPORT_251_addr = 8'hfb;
  assign ram_3_MPORT_251_mask = 1'h1;
  assign ram_3_MPORT_251_en = reset;
  assign ram_3_MPORT_252_data = 2'h0;
  assign ram_3_MPORT_252_addr = 8'hfc;
  assign ram_3_MPORT_252_mask = 1'h1;
  assign ram_3_MPORT_252_en = reset;
  assign ram_3_MPORT_253_data = 2'h0;
  assign ram_3_MPORT_253_addr = 8'hfd;
  assign ram_3_MPORT_253_mask = 1'h1;
  assign ram_3_MPORT_253_en = reset;
  assign ram_3_MPORT_254_data = 2'h0;
  assign ram_3_MPORT_254_addr = 8'hfe;
  assign ram_3_MPORT_254_mask = 1'h1;
  assign ram_3_MPORT_254_en = reset;
  assign ram_3_MPORT_255_data = 2'h0;
  assign ram_3_MPORT_255_addr = 8'hff;
  assign ram_3_MPORT_255_mask = 1'h1;
  assign ram_3_MPORT_255_en = reset;
  assign ram_3_MPORT_256_data = io_wdata[7:6];
  assign ram_3_MPORT_256_addr = io_addr;
  assign ram_3_MPORT_256_mask = io_wmask[3];
  assign ram_3_MPORT_256_en = io_rw;
  assign io_rdata = {io_rdata_hi,io_rdata_lo}; // @[SRAM.scala 75:39]
  always @(posedge clock) begin
    if (ram_0_MPORT_en & ram_0_MPORT_mask) begin
      ram_0[ram_0_MPORT_addr] <= ram_0_MPORT_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_1_en & ram_0_MPORT_1_mask) begin
      ram_0[ram_0_MPORT_1_addr] <= ram_0_MPORT_1_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_2_en & ram_0_MPORT_2_mask) begin
      ram_0[ram_0_MPORT_2_addr] <= ram_0_MPORT_2_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_3_en & ram_0_MPORT_3_mask) begin
      ram_0[ram_0_MPORT_3_addr] <= ram_0_MPORT_3_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_4_en & ram_0_MPORT_4_mask) begin
      ram_0[ram_0_MPORT_4_addr] <= ram_0_MPORT_4_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_5_en & ram_0_MPORT_5_mask) begin
      ram_0[ram_0_MPORT_5_addr] <= ram_0_MPORT_5_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_6_en & ram_0_MPORT_6_mask) begin
      ram_0[ram_0_MPORT_6_addr] <= ram_0_MPORT_6_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_7_en & ram_0_MPORT_7_mask) begin
      ram_0[ram_0_MPORT_7_addr] <= ram_0_MPORT_7_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_8_en & ram_0_MPORT_8_mask) begin
      ram_0[ram_0_MPORT_8_addr] <= ram_0_MPORT_8_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_9_en & ram_0_MPORT_9_mask) begin
      ram_0[ram_0_MPORT_9_addr] <= ram_0_MPORT_9_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_10_en & ram_0_MPORT_10_mask) begin
      ram_0[ram_0_MPORT_10_addr] <= ram_0_MPORT_10_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_11_en & ram_0_MPORT_11_mask) begin
      ram_0[ram_0_MPORT_11_addr] <= ram_0_MPORT_11_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_12_en & ram_0_MPORT_12_mask) begin
      ram_0[ram_0_MPORT_12_addr] <= ram_0_MPORT_12_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_13_en & ram_0_MPORT_13_mask) begin
      ram_0[ram_0_MPORT_13_addr] <= ram_0_MPORT_13_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_14_en & ram_0_MPORT_14_mask) begin
      ram_0[ram_0_MPORT_14_addr] <= ram_0_MPORT_14_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_15_en & ram_0_MPORT_15_mask) begin
      ram_0[ram_0_MPORT_15_addr] <= ram_0_MPORT_15_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_16_en & ram_0_MPORT_16_mask) begin
      ram_0[ram_0_MPORT_16_addr] <= ram_0_MPORT_16_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_17_en & ram_0_MPORT_17_mask) begin
      ram_0[ram_0_MPORT_17_addr] <= ram_0_MPORT_17_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_18_en & ram_0_MPORT_18_mask) begin
      ram_0[ram_0_MPORT_18_addr] <= ram_0_MPORT_18_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_19_en & ram_0_MPORT_19_mask) begin
      ram_0[ram_0_MPORT_19_addr] <= ram_0_MPORT_19_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_20_en & ram_0_MPORT_20_mask) begin
      ram_0[ram_0_MPORT_20_addr] <= ram_0_MPORT_20_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_21_en & ram_0_MPORT_21_mask) begin
      ram_0[ram_0_MPORT_21_addr] <= ram_0_MPORT_21_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_22_en & ram_0_MPORT_22_mask) begin
      ram_0[ram_0_MPORT_22_addr] <= ram_0_MPORT_22_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_23_en & ram_0_MPORT_23_mask) begin
      ram_0[ram_0_MPORT_23_addr] <= ram_0_MPORT_23_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_24_en & ram_0_MPORT_24_mask) begin
      ram_0[ram_0_MPORT_24_addr] <= ram_0_MPORT_24_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_25_en & ram_0_MPORT_25_mask) begin
      ram_0[ram_0_MPORT_25_addr] <= ram_0_MPORT_25_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_26_en & ram_0_MPORT_26_mask) begin
      ram_0[ram_0_MPORT_26_addr] <= ram_0_MPORT_26_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_27_en & ram_0_MPORT_27_mask) begin
      ram_0[ram_0_MPORT_27_addr] <= ram_0_MPORT_27_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_28_en & ram_0_MPORT_28_mask) begin
      ram_0[ram_0_MPORT_28_addr] <= ram_0_MPORT_28_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_29_en & ram_0_MPORT_29_mask) begin
      ram_0[ram_0_MPORT_29_addr] <= ram_0_MPORT_29_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_30_en & ram_0_MPORT_30_mask) begin
      ram_0[ram_0_MPORT_30_addr] <= ram_0_MPORT_30_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_31_en & ram_0_MPORT_31_mask) begin
      ram_0[ram_0_MPORT_31_addr] <= ram_0_MPORT_31_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_32_en & ram_0_MPORT_32_mask) begin
      ram_0[ram_0_MPORT_32_addr] <= ram_0_MPORT_32_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_33_en & ram_0_MPORT_33_mask) begin
      ram_0[ram_0_MPORT_33_addr] <= ram_0_MPORT_33_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_34_en & ram_0_MPORT_34_mask) begin
      ram_0[ram_0_MPORT_34_addr] <= ram_0_MPORT_34_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_35_en & ram_0_MPORT_35_mask) begin
      ram_0[ram_0_MPORT_35_addr] <= ram_0_MPORT_35_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_36_en & ram_0_MPORT_36_mask) begin
      ram_0[ram_0_MPORT_36_addr] <= ram_0_MPORT_36_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_37_en & ram_0_MPORT_37_mask) begin
      ram_0[ram_0_MPORT_37_addr] <= ram_0_MPORT_37_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_38_en & ram_0_MPORT_38_mask) begin
      ram_0[ram_0_MPORT_38_addr] <= ram_0_MPORT_38_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_39_en & ram_0_MPORT_39_mask) begin
      ram_0[ram_0_MPORT_39_addr] <= ram_0_MPORT_39_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_40_en & ram_0_MPORT_40_mask) begin
      ram_0[ram_0_MPORT_40_addr] <= ram_0_MPORT_40_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_41_en & ram_0_MPORT_41_mask) begin
      ram_0[ram_0_MPORT_41_addr] <= ram_0_MPORT_41_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_42_en & ram_0_MPORT_42_mask) begin
      ram_0[ram_0_MPORT_42_addr] <= ram_0_MPORT_42_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_43_en & ram_0_MPORT_43_mask) begin
      ram_0[ram_0_MPORT_43_addr] <= ram_0_MPORT_43_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_44_en & ram_0_MPORT_44_mask) begin
      ram_0[ram_0_MPORT_44_addr] <= ram_0_MPORT_44_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_45_en & ram_0_MPORT_45_mask) begin
      ram_0[ram_0_MPORT_45_addr] <= ram_0_MPORT_45_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_46_en & ram_0_MPORT_46_mask) begin
      ram_0[ram_0_MPORT_46_addr] <= ram_0_MPORT_46_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_47_en & ram_0_MPORT_47_mask) begin
      ram_0[ram_0_MPORT_47_addr] <= ram_0_MPORT_47_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_48_en & ram_0_MPORT_48_mask) begin
      ram_0[ram_0_MPORT_48_addr] <= ram_0_MPORT_48_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_49_en & ram_0_MPORT_49_mask) begin
      ram_0[ram_0_MPORT_49_addr] <= ram_0_MPORT_49_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_50_en & ram_0_MPORT_50_mask) begin
      ram_0[ram_0_MPORT_50_addr] <= ram_0_MPORT_50_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_51_en & ram_0_MPORT_51_mask) begin
      ram_0[ram_0_MPORT_51_addr] <= ram_0_MPORT_51_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_52_en & ram_0_MPORT_52_mask) begin
      ram_0[ram_0_MPORT_52_addr] <= ram_0_MPORT_52_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_53_en & ram_0_MPORT_53_mask) begin
      ram_0[ram_0_MPORT_53_addr] <= ram_0_MPORT_53_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_54_en & ram_0_MPORT_54_mask) begin
      ram_0[ram_0_MPORT_54_addr] <= ram_0_MPORT_54_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_55_en & ram_0_MPORT_55_mask) begin
      ram_0[ram_0_MPORT_55_addr] <= ram_0_MPORT_55_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_56_en & ram_0_MPORT_56_mask) begin
      ram_0[ram_0_MPORT_56_addr] <= ram_0_MPORT_56_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_57_en & ram_0_MPORT_57_mask) begin
      ram_0[ram_0_MPORT_57_addr] <= ram_0_MPORT_57_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_58_en & ram_0_MPORT_58_mask) begin
      ram_0[ram_0_MPORT_58_addr] <= ram_0_MPORT_58_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_59_en & ram_0_MPORT_59_mask) begin
      ram_0[ram_0_MPORT_59_addr] <= ram_0_MPORT_59_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_60_en & ram_0_MPORT_60_mask) begin
      ram_0[ram_0_MPORT_60_addr] <= ram_0_MPORT_60_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_61_en & ram_0_MPORT_61_mask) begin
      ram_0[ram_0_MPORT_61_addr] <= ram_0_MPORT_61_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_62_en & ram_0_MPORT_62_mask) begin
      ram_0[ram_0_MPORT_62_addr] <= ram_0_MPORT_62_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_63_en & ram_0_MPORT_63_mask) begin
      ram_0[ram_0_MPORT_63_addr] <= ram_0_MPORT_63_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_64_en & ram_0_MPORT_64_mask) begin
      ram_0[ram_0_MPORT_64_addr] <= ram_0_MPORT_64_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_65_en & ram_0_MPORT_65_mask) begin
      ram_0[ram_0_MPORT_65_addr] <= ram_0_MPORT_65_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_66_en & ram_0_MPORT_66_mask) begin
      ram_0[ram_0_MPORT_66_addr] <= ram_0_MPORT_66_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_67_en & ram_0_MPORT_67_mask) begin
      ram_0[ram_0_MPORT_67_addr] <= ram_0_MPORT_67_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_68_en & ram_0_MPORT_68_mask) begin
      ram_0[ram_0_MPORT_68_addr] <= ram_0_MPORT_68_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_69_en & ram_0_MPORT_69_mask) begin
      ram_0[ram_0_MPORT_69_addr] <= ram_0_MPORT_69_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_70_en & ram_0_MPORT_70_mask) begin
      ram_0[ram_0_MPORT_70_addr] <= ram_0_MPORT_70_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_71_en & ram_0_MPORT_71_mask) begin
      ram_0[ram_0_MPORT_71_addr] <= ram_0_MPORT_71_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_72_en & ram_0_MPORT_72_mask) begin
      ram_0[ram_0_MPORT_72_addr] <= ram_0_MPORT_72_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_73_en & ram_0_MPORT_73_mask) begin
      ram_0[ram_0_MPORT_73_addr] <= ram_0_MPORT_73_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_74_en & ram_0_MPORT_74_mask) begin
      ram_0[ram_0_MPORT_74_addr] <= ram_0_MPORT_74_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_75_en & ram_0_MPORT_75_mask) begin
      ram_0[ram_0_MPORT_75_addr] <= ram_0_MPORT_75_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_76_en & ram_0_MPORT_76_mask) begin
      ram_0[ram_0_MPORT_76_addr] <= ram_0_MPORT_76_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_77_en & ram_0_MPORT_77_mask) begin
      ram_0[ram_0_MPORT_77_addr] <= ram_0_MPORT_77_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_78_en & ram_0_MPORT_78_mask) begin
      ram_0[ram_0_MPORT_78_addr] <= ram_0_MPORT_78_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_79_en & ram_0_MPORT_79_mask) begin
      ram_0[ram_0_MPORT_79_addr] <= ram_0_MPORT_79_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_80_en & ram_0_MPORT_80_mask) begin
      ram_0[ram_0_MPORT_80_addr] <= ram_0_MPORT_80_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_81_en & ram_0_MPORT_81_mask) begin
      ram_0[ram_0_MPORT_81_addr] <= ram_0_MPORT_81_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_82_en & ram_0_MPORT_82_mask) begin
      ram_0[ram_0_MPORT_82_addr] <= ram_0_MPORT_82_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_83_en & ram_0_MPORT_83_mask) begin
      ram_0[ram_0_MPORT_83_addr] <= ram_0_MPORT_83_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_84_en & ram_0_MPORT_84_mask) begin
      ram_0[ram_0_MPORT_84_addr] <= ram_0_MPORT_84_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_85_en & ram_0_MPORT_85_mask) begin
      ram_0[ram_0_MPORT_85_addr] <= ram_0_MPORT_85_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_86_en & ram_0_MPORT_86_mask) begin
      ram_0[ram_0_MPORT_86_addr] <= ram_0_MPORT_86_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_87_en & ram_0_MPORT_87_mask) begin
      ram_0[ram_0_MPORT_87_addr] <= ram_0_MPORT_87_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_88_en & ram_0_MPORT_88_mask) begin
      ram_0[ram_0_MPORT_88_addr] <= ram_0_MPORT_88_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_89_en & ram_0_MPORT_89_mask) begin
      ram_0[ram_0_MPORT_89_addr] <= ram_0_MPORT_89_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_90_en & ram_0_MPORT_90_mask) begin
      ram_0[ram_0_MPORT_90_addr] <= ram_0_MPORT_90_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_91_en & ram_0_MPORT_91_mask) begin
      ram_0[ram_0_MPORT_91_addr] <= ram_0_MPORT_91_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_92_en & ram_0_MPORT_92_mask) begin
      ram_0[ram_0_MPORT_92_addr] <= ram_0_MPORT_92_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_93_en & ram_0_MPORT_93_mask) begin
      ram_0[ram_0_MPORT_93_addr] <= ram_0_MPORT_93_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_94_en & ram_0_MPORT_94_mask) begin
      ram_0[ram_0_MPORT_94_addr] <= ram_0_MPORT_94_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_95_en & ram_0_MPORT_95_mask) begin
      ram_0[ram_0_MPORT_95_addr] <= ram_0_MPORT_95_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_96_en & ram_0_MPORT_96_mask) begin
      ram_0[ram_0_MPORT_96_addr] <= ram_0_MPORT_96_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_97_en & ram_0_MPORT_97_mask) begin
      ram_0[ram_0_MPORT_97_addr] <= ram_0_MPORT_97_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_98_en & ram_0_MPORT_98_mask) begin
      ram_0[ram_0_MPORT_98_addr] <= ram_0_MPORT_98_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_99_en & ram_0_MPORT_99_mask) begin
      ram_0[ram_0_MPORT_99_addr] <= ram_0_MPORT_99_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_100_en & ram_0_MPORT_100_mask) begin
      ram_0[ram_0_MPORT_100_addr] <= ram_0_MPORT_100_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_101_en & ram_0_MPORT_101_mask) begin
      ram_0[ram_0_MPORT_101_addr] <= ram_0_MPORT_101_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_102_en & ram_0_MPORT_102_mask) begin
      ram_0[ram_0_MPORT_102_addr] <= ram_0_MPORT_102_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_103_en & ram_0_MPORT_103_mask) begin
      ram_0[ram_0_MPORT_103_addr] <= ram_0_MPORT_103_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_104_en & ram_0_MPORT_104_mask) begin
      ram_0[ram_0_MPORT_104_addr] <= ram_0_MPORT_104_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_105_en & ram_0_MPORT_105_mask) begin
      ram_0[ram_0_MPORT_105_addr] <= ram_0_MPORT_105_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_106_en & ram_0_MPORT_106_mask) begin
      ram_0[ram_0_MPORT_106_addr] <= ram_0_MPORT_106_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_107_en & ram_0_MPORT_107_mask) begin
      ram_0[ram_0_MPORT_107_addr] <= ram_0_MPORT_107_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_108_en & ram_0_MPORT_108_mask) begin
      ram_0[ram_0_MPORT_108_addr] <= ram_0_MPORT_108_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_109_en & ram_0_MPORT_109_mask) begin
      ram_0[ram_0_MPORT_109_addr] <= ram_0_MPORT_109_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_110_en & ram_0_MPORT_110_mask) begin
      ram_0[ram_0_MPORT_110_addr] <= ram_0_MPORT_110_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_111_en & ram_0_MPORT_111_mask) begin
      ram_0[ram_0_MPORT_111_addr] <= ram_0_MPORT_111_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_112_en & ram_0_MPORT_112_mask) begin
      ram_0[ram_0_MPORT_112_addr] <= ram_0_MPORT_112_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_113_en & ram_0_MPORT_113_mask) begin
      ram_0[ram_0_MPORT_113_addr] <= ram_0_MPORT_113_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_114_en & ram_0_MPORT_114_mask) begin
      ram_0[ram_0_MPORT_114_addr] <= ram_0_MPORT_114_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_115_en & ram_0_MPORT_115_mask) begin
      ram_0[ram_0_MPORT_115_addr] <= ram_0_MPORT_115_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_116_en & ram_0_MPORT_116_mask) begin
      ram_0[ram_0_MPORT_116_addr] <= ram_0_MPORT_116_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_117_en & ram_0_MPORT_117_mask) begin
      ram_0[ram_0_MPORT_117_addr] <= ram_0_MPORT_117_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_118_en & ram_0_MPORT_118_mask) begin
      ram_0[ram_0_MPORT_118_addr] <= ram_0_MPORT_118_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_119_en & ram_0_MPORT_119_mask) begin
      ram_0[ram_0_MPORT_119_addr] <= ram_0_MPORT_119_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_120_en & ram_0_MPORT_120_mask) begin
      ram_0[ram_0_MPORT_120_addr] <= ram_0_MPORT_120_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_121_en & ram_0_MPORT_121_mask) begin
      ram_0[ram_0_MPORT_121_addr] <= ram_0_MPORT_121_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_122_en & ram_0_MPORT_122_mask) begin
      ram_0[ram_0_MPORT_122_addr] <= ram_0_MPORT_122_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_123_en & ram_0_MPORT_123_mask) begin
      ram_0[ram_0_MPORT_123_addr] <= ram_0_MPORT_123_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_124_en & ram_0_MPORT_124_mask) begin
      ram_0[ram_0_MPORT_124_addr] <= ram_0_MPORT_124_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_125_en & ram_0_MPORT_125_mask) begin
      ram_0[ram_0_MPORT_125_addr] <= ram_0_MPORT_125_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_126_en & ram_0_MPORT_126_mask) begin
      ram_0[ram_0_MPORT_126_addr] <= ram_0_MPORT_126_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_127_en & ram_0_MPORT_127_mask) begin
      ram_0[ram_0_MPORT_127_addr] <= ram_0_MPORT_127_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_128_en & ram_0_MPORT_128_mask) begin
      ram_0[ram_0_MPORT_128_addr] <= ram_0_MPORT_128_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_129_en & ram_0_MPORT_129_mask) begin
      ram_0[ram_0_MPORT_129_addr] <= ram_0_MPORT_129_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_130_en & ram_0_MPORT_130_mask) begin
      ram_0[ram_0_MPORT_130_addr] <= ram_0_MPORT_130_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_131_en & ram_0_MPORT_131_mask) begin
      ram_0[ram_0_MPORT_131_addr] <= ram_0_MPORT_131_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_132_en & ram_0_MPORT_132_mask) begin
      ram_0[ram_0_MPORT_132_addr] <= ram_0_MPORT_132_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_133_en & ram_0_MPORT_133_mask) begin
      ram_0[ram_0_MPORT_133_addr] <= ram_0_MPORT_133_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_134_en & ram_0_MPORT_134_mask) begin
      ram_0[ram_0_MPORT_134_addr] <= ram_0_MPORT_134_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_135_en & ram_0_MPORT_135_mask) begin
      ram_0[ram_0_MPORT_135_addr] <= ram_0_MPORT_135_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_136_en & ram_0_MPORT_136_mask) begin
      ram_0[ram_0_MPORT_136_addr] <= ram_0_MPORT_136_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_137_en & ram_0_MPORT_137_mask) begin
      ram_0[ram_0_MPORT_137_addr] <= ram_0_MPORT_137_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_138_en & ram_0_MPORT_138_mask) begin
      ram_0[ram_0_MPORT_138_addr] <= ram_0_MPORT_138_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_139_en & ram_0_MPORT_139_mask) begin
      ram_0[ram_0_MPORT_139_addr] <= ram_0_MPORT_139_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_140_en & ram_0_MPORT_140_mask) begin
      ram_0[ram_0_MPORT_140_addr] <= ram_0_MPORT_140_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_141_en & ram_0_MPORT_141_mask) begin
      ram_0[ram_0_MPORT_141_addr] <= ram_0_MPORT_141_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_142_en & ram_0_MPORT_142_mask) begin
      ram_0[ram_0_MPORT_142_addr] <= ram_0_MPORT_142_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_143_en & ram_0_MPORT_143_mask) begin
      ram_0[ram_0_MPORT_143_addr] <= ram_0_MPORT_143_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_144_en & ram_0_MPORT_144_mask) begin
      ram_0[ram_0_MPORT_144_addr] <= ram_0_MPORT_144_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_145_en & ram_0_MPORT_145_mask) begin
      ram_0[ram_0_MPORT_145_addr] <= ram_0_MPORT_145_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_146_en & ram_0_MPORT_146_mask) begin
      ram_0[ram_0_MPORT_146_addr] <= ram_0_MPORT_146_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_147_en & ram_0_MPORT_147_mask) begin
      ram_0[ram_0_MPORT_147_addr] <= ram_0_MPORT_147_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_148_en & ram_0_MPORT_148_mask) begin
      ram_0[ram_0_MPORT_148_addr] <= ram_0_MPORT_148_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_149_en & ram_0_MPORT_149_mask) begin
      ram_0[ram_0_MPORT_149_addr] <= ram_0_MPORT_149_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_150_en & ram_0_MPORT_150_mask) begin
      ram_0[ram_0_MPORT_150_addr] <= ram_0_MPORT_150_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_151_en & ram_0_MPORT_151_mask) begin
      ram_0[ram_0_MPORT_151_addr] <= ram_0_MPORT_151_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_152_en & ram_0_MPORT_152_mask) begin
      ram_0[ram_0_MPORT_152_addr] <= ram_0_MPORT_152_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_153_en & ram_0_MPORT_153_mask) begin
      ram_0[ram_0_MPORT_153_addr] <= ram_0_MPORT_153_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_154_en & ram_0_MPORT_154_mask) begin
      ram_0[ram_0_MPORT_154_addr] <= ram_0_MPORT_154_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_155_en & ram_0_MPORT_155_mask) begin
      ram_0[ram_0_MPORT_155_addr] <= ram_0_MPORT_155_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_156_en & ram_0_MPORT_156_mask) begin
      ram_0[ram_0_MPORT_156_addr] <= ram_0_MPORT_156_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_157_en & ram_0_MPORT_157_mask) begin
      ram_0[ram_0_MPORT_157_addr] <= ram_0_MPORT_157_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_158_en & ram_0_MPORT_158_mask) begin
      ram_0[ram_0_MPORT_158_addr] <= ram_0_MPORT_158_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_159_en & ram_0_MPORT_159_mask) begin
      ram_0[ram_0_MPORT_159_addr] <= ram_0_MPORT_159_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_160_en & ram_0_MPORT_160_mask) begin
      ram_0[ram_0_MPORT_160_addr] <= ram_0_MPORT_160_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_161_en & ram_0_MPORT_161_mask) begin
      ram_0[ram_0_MPORT_161_addr] <= ram_0_MPORT_161_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_162_en & ram_0_MPORT_162_mask) begin
      ram_0[ram_0_MPORT_162_addr] <= ram_0_MPORT_162_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_163_en & ram_0_MPORT_163_mask) begin
      ram_0[ram_0_MPORT_163_addr] <= ram_0_MPORT_163_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_164_en & ram_0_MPORT_164_mask) begin
      ram_0[ram_0_MPORT_164_addr] <= ram_0_MPORT_164_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_165_en & ram_0_MPORT_165_mask) begin
      ram_0[ram_0_MPORT_165_addr] <= ram_0_MPORT_165_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_166_en & ram_0_MPORT_166_mask) begin
      ram_0[ram_0_MPORT_166_addr] <= ram_0_MPORT_166_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_167_en & ram_0_MPORT_167_mask) begin
      ram_0[ram_0_MPORT_167_addr] <= ram_0_MPORT_167_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_168_en & ram_0_MPORT_168_mask) begin
      ram_0[ram_0_MPORT_168_addr] <= ram_0_MPORT_168_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_169_en & ram_0_MPORT_169_mask) begin
      ram_0[ram_0_MPORT_169_addr] <= ram_0_MPORT_169_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_170_en & ram_0_MPORT_170_mask) begin
      ram_0[ram_0_MPORT_170_addr] <= ram_0_MPORT_170_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_171_en & ram_0_MPORT_171_mask) begin
      ram_0[ram_0_MPORT_171_addr] <= ram_0_MPORT_171_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_172_en & ram_0_MPORT_172_mask) begin
      ram_0[ram_0_MPORT_172_addr] <= ram_0_MPORT_172_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_173_en & ram_0_MPORT_173_mask) begin
      ram_0[ram_0_MPORT_173_addr] <= ram_0_MPORT_173_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_174_en & ram_0_MPORT_174_mask) begin
      ram_0[ram_0_MPORT_174_addr] <= ram_0_MPORT_174_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_175_en & ram_0_MPORT_175_mask) begin
      ram_0[ram_0_MPORT_175_addr] <= ram_0_MPORT_175_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_176_en & ram_0_MPORT_176_mask) begin
      ram_0[ram_0_MPORT_176_addr] <= ram_0_MPORT_176_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_177_en & ram_0_MPORT_177_mask) begin
      ram_0[ram_0_MPORT_177_addr] <= ram_0_MPORT_177_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_178_en & ram_0_MPORT_178_mask) begin
      ram_0[ram_0_MPORT_178_addr] <= ram_0_MPORT_178_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_179_en & ram_0_MPORT_179_mask) begin
      ram_0[ram_0_MPORT_179_addr] <= ram_0_MPORT_179_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_180_en & ram_0_MPORT_180_mask) begin
      ram_0[ram_0_MPORT_180_addr] <= ram_0_MPORT_180_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_181_en & ram_0_MPORT_181_mask) begin
      ram_0[ram_0_MPORT_181_addr] <= ram_0_MPORT_181_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_182_en & ram_0_MPORT_182_mask) begin
      ram_0[ram_0_MPORT_182_addr] <= ram_0_MPORT_182_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_183_en & ram_0_MPORT_183_mask) begin
      ram_0[ram_0_MPORT_183_addr] <= ram_0_MPORT_183_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_184_en & ram_0_MPORT_184_mask) begin
      ram_0[ram_0_MPORT_184_addr] <= ram_0_MPORT_184_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_185_en & ram_0_MPORT_185_mask) begin
      ram_0[ram_0_MPORT_185_addr] <= ram_0_MPORT_185_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_186_en & ram_0_MPORT_186_mask) begin
      ram_0[ram_0_MPORT_186_addr] <= ram_0_MPORT_186_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_187_en & ram_0_MPORT_187_mask) begin
      ram_0[ram_0_MPORT_187_addr] <= ram_0_MPORT_187_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_188_en & ram_0_MPORT_188_mask) begin
      ram_0[ram_0_MPORT_188_addr] <= ram_0_MPORT_188_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_189_en & ram_0_MPORT_189_mask) begin
      ram_0[ram_0_MPORT_189_addr] <= ram_0_MPORT_189_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_190_en & ram_0_MPORT_190_mask) begin
      ram_0[ram_0_MPORT_190_addr] <= ram_0_MPORT_190_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_191_en & ram_0_MPORT_191_mask) begin
      ram_0[ram_0_MPORT_191_addr] <= ram_0_MPORT_191_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_192_en & ram_0_MPORT_192_mask) begin
      ram_0[ram_0_MPORT_192_addr] <= ram_0_MPORT_192_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_193_en & ram_0_MPORT_193_mask) begin
      ram_0[ram_0_MPORT_193_addr] <= ram_0_MPORT_193_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_194_en & ram_0_MPORT_194_mask) begin
      ram_0[ram_0_MPORT_194_addr] <= ram_0_MPORT_194_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_195_en & ram_0_MPORT_195_mask) begin
      ram_0[ram_0_MPORT_195_addr] <= ram_0_MPORT_195_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_196_en & ram_0_MPORT_196_mask) begin
      ram_0[ram_0_MPORT_196_addr] <= ram_0_MPORT_196_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_197_en & ram_0_MPORT_197_mask) begin
      ram_0[ram_0_MPORT_197_addr] <= ram_0_MPORT_197_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_198_en & ram_0_MPORT_198_mask) begin
      ram_0[ram_0_MPORT_198_addr] <= ram_0_MPORT_198_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_199_en & ram_0_MPORT_199_mask) begin
      ram_0[ram_0_MPORT_199_addr] <= ram_0_MPORT_199_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_200_en & ram_0_MPORT_200_mask) begin
      ram_0[ram_0_MPORT_200_addr] <= ram_0_MPORT_200_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_201_en & ram_0_MPORT_201_mask) begin
      ram_0[ram_0_MPORT_201_addr] <= ram_0_MPORT_201_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_202_en & ram_0_MPORT_202_mask) begin
      ram_0[ram_0_MPORT_202_addr] <= ram_0_MPORT_202_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_203_en & ram_0_MPORT_203_mask) begin
      ram_0[ram_0_MPORT_203_addr] <= ram_0_MPORT_203_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_204_en & ram_0_MPORT_204_mask) begin
      ram_0[ram_0_MPORT_204_addr] <= ram_0_MPORT_204_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_205_en & ram_0_MPORT_205_mask) begin
      ram_0[ram_0_MPORT_205_addr] <= ram_0_MPORT_205_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_206_en & ram_0_MPORT_206_mask) begin
      ram_0[ram_0_MPORT_206_addr] <= ram_0_MPORT_206_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_207_en & ram_0_MPORT_207_mask) begin
      ram_0[ram_0_MPORT_207_addr] <= ram_0_MPORT_207_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_208_en & ram_0_MPORT_208_mask) begin
      ram_0[ram_0_MPORT_208_addr] <= ram_0_MPORT_208_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_209_en & ram_0_MPORT_209_mask) begin
      ram_0[ram_0_MPORT_209_addr] <= ram_0_MPORT_209_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_210_en & ram_0_MPORT_210_mask) begin
      ram_0[ram_0_MPORT_210_addr] <= ram_0_MPORT_210_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_211_en & ram_0_MPORT_211_mask) begin
      ram_0[ram_0_MPORT_211_addr] <= ram_0_MPORT_211_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_212_en & ram_0_MPORT_212_mask) begin
      ram_0[ram_0_MPORT_212_addr] <= ram_0_MPORT_212_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_213_en & ram_0_MPORT_213_mask) begin
      ram_0[ram_0_MPORT_213_addr] <= ram_0_MPORT_213_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_214_en & ram_0_MPORT_214_mask) begin
      ram_0[ram_0_MPORT_214_addr] <= ram_0_MPORT_214_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_215_en & ram_0_MPORT_215_mask) begin
      ram_0[ram_0_MPORT_215_addr] <= ram_0_MPORT_215_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_216_en & ram_0_MPORT_216_mask) begin
      ram_0[ram_0_MPORT_216_addr] <= ram_0_MPORT_216_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_217_en & ram_0_MPORT_217_mask) begin
      ram_0[ram_0_MPORT_217_addr] <= ram_0_MPORT_217_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_218_en & ram_0_MPORT_218_mask) begin
      ram_0[ram_0_MPORT_218_addr] <= ram_0_MPORT_218_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_219_en & ram_0_MPORT_219_mask) begin
      ram_0[ram_0_MPORT_219_addr] <= ram_0_MPORT_219_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_220_en & ram_0_MPORT_220_mask) begin
      ram_0[ram_0_MPORT_220_addr] <= ram_0_MPORT_220_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_221_en & ram_0_MPORT_221_mask) begin
      ram_0[ram_0_MPORT_221_addr] <= ram_0_MPORT_221_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_222_en & ram_0_MPORT_222_mask) begin
      ram_0[ram_0_MPORT_222_addr] <= ram_0_MPORT_222_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_223_en & ram_0_MPORT_223_mask) begin
      ram_0[ram_0_MPORT_223_addr] <= ram_0_MPORT_223_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_224_en & ram_0_MPORT_224_mask) begin
      ram_0[ram_0_MPORT_224_addr] <= ram_0_MPORT_224_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_225_en & ram_0_MPORT_225_mask) begin
      ram_0[ram_0_MPORT_225_addr] <= ram_0_MPORT_225_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_226_en & ram_0_MPORT_226_mask) begin
      ram_0[ram_0_MPORT_226_addr] <= ram_0_MPORT_226_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_227_en & ram_0_MPORT_227_mask) begin
      ram_0[ram_0_MPORT_227_addr] <= ram_0_MPORT_227_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_228_en & ram_0_MPORT_228_mask) begin
      ram_0[ram_0_MPORT_228_addr] <= ram_0_MPORT_228_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_229_en & ram_0_MPORT_229_mask) begin
      ram_0[ram_0_MPORT_229_addr] <= ram_0_MPORT_229_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_230_en & ram_0_MPORT_230_mask) begin
      ram_0[ram_0_MPORT_230_addr] <= ram_0_MPORT_230_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_231_en & ram_0_MPORT_231_mask) begin
      ram_0[ram_0_MPORT_231_addr] <= ram_0_MPORT_231_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_232_en & ram_0_MPORT_232_mask) begin
      ram_0[ram_0_MPORT_232_addr] <= ram_0_MPORT_232_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_233_en & ram_0_MPORT_233_mask) begin
      ram_0[ram_0_MPORT_233_addr] <= ram_0_MPORT_233_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_234_en & ram_0_MPORT_234_mask) begin
      ram_0[ram_0_MPORT_234_addr] <= ram_0_MPORT_234_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_235_en & ram_0_MPORT_235_mask) begin
      ram_0[ram_0_MPORT_235_addr] <= ram_0_MPORT_235_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_236_en & ram_0_MPORT_236_mask) begin
      ram_0[ram_0_MPORT_236_addr] <= ram_0_MPORT_236_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_237_en & ram_0_MPORT_237_mask) begin
      ram_0[ram_0_MPORT_237_addr] <= ram_0_MPORT_237_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_238_en & ram_0_MPORT_238_mask) begin
      ram_0[ram_0_MPORT_238_addr] <= ram_0_MPORT_238_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_239_en & ram_0_MPORT_239_mask) begin
      ram_0[ram_0_MPORT_239_addr] <= ram_0_MPORT_239_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_240_en & ram_0_MPORT_240_mask) begin
      ram_0[ram_0_MPORT_240_addr] <= ram_0_MPORT_240_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_241_en & ram_0_MPORT_241_mask) begin
      ram_0[ram_0_MPORT_241_addr] <= ram_0_MPORT_241_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_242_en & ram_0_MPORT_242_mask) begin
      ram_0[ram_0_MPORT_242_addr] <= ram_0_MPORT_242_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_243_en & ram_0_MPORT_243_mask) begin
      ram_0[ram_0_MPORT_243_addr] <= ram_0_MPORT_243_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_244_en & ram_0_MPORT_244_mask) begin
      ram_0[ram_0_MPORT_244_addr] <= ram_0_MPORT_244_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_245_en & ram_0_MPORT_245_mask) begin
      ram_0[ram_0_MPORT_245_addr] <= ram_0_MPORT_245_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_246_en & ram_0_MPORT_246_mask) begin
      ram_0[ram_0_MPORT_246_addr] <= ram_0_MPORT_246_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_247_en & ram_0_MPORT_247_mask) begin
      ram_0[ram_0_MPORT_247_addr] <= ram_0_MPORT_247_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_248_en & ram_0_MPORT_248_mask) begin
      ram_0[ram_0_MPORT_248_addr] <= ram_0_MPORT_248_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_249_en & ram_0_MPORT_249_mask) begin
      ram_0[ram_0_MPORT_249_addr] <= ram_0_MPORT_249_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_250_en & ram_0_MPORT_250_mask) begin
      ram_0[ram_0_MPORT_250_addr] <= ram_0_MPORT_250_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_251_en & ram_0_MPORT_251_mask) begin
      ram_0[ram_0_MPORT_251_addr] <= ram_0_MPORT_251_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_252_en & ram_0_MPORT_252_mask) begin
      ram_0[ram_0_MPORT_252_addr] <= ram_0_MPORT_252_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_253_en & ram_0_MPORT_253_mask) begin
      ram_0[ram_0_MPORT_253_addr] <= ram_0_MPORT_253_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_254_en & ram_0_MPORT_254_mask) begin
      ram_0[ram_0_MPORT_254_addr] <= ram_0_MPORT_254_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_255_en & ram_0_MPORT_255_mask) begin
      ram_0[ram_0_MPORT_255_addr] <= ram_0_MPORT_255_data; // @[SRAM.scala 36:26]
    end
    if (ram_0_MPORT_256_en & ram_0_MPORT_256_mask) begin
      ram_0[ram_0_MPORT_256_addr] <= ram_0_MPORT_256_data; // @[SRAM.scala 36:26]
    end
    if (io_rw) begin
      ram_0_io_rdata_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      ram_0_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    end
    if (io_rw ? 1'h0 : 1'h1) begin
      ram_0_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
    if (ram_1_MPORT_en & ram_1_MPORT_mask) begin
      ram_1[ram_1_MPORT_addr] <= ram_1_MPORT_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_1_en & ram_1_MPORT_1_mask) begin
      ram_1[ram_1_MPORT_1_addr] <= ram_1_MPORT_1_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_2_en & ram_1_MPORT_2_mask) begin
      ram_1[ram_1_MPORT_2_addr] <= ram_1_MPORT_2_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_3_en & ram_1_MPORT_3_mask) begin
      ram_1[ram_1_MPORT_3_addr] <= ram_1_MPORT_3_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_4_en & ram_1_MPORT_4_mask) begin
      ram_1[ram_1_MPORT_4_addr] <= ram_1_MPORT_4_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_5_en & ram_1_MPORT_5_mask) begin
      ram_1[ram_1_MPORT_5_addr] <= ram_1_MPORT_5_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_6_en & ram_1_MPORT_6_mask) begin
      ram_1[ram_1_MPORT_6_addr] <= ram_1_MPORT_6_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_7_en & ram_1_MPORT_7_mask) begin
      ram_1[ram_1_MPORT_7_addr] <= ram_1_MPORT_7_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_8_en & ram_1_MPORT_8_mask) begin
      ram_1[ram_1_MPORT_8_addr] <= ram_1_MPORT_8_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_9_en & ram_1_MPORT_9_mask) begin
      ram_1[ram_1_MPORT_9_addr] <= ram_1_MPORT_9_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_10_en & ram_1_MPORT_10_mask) begin
      ram_1[ram_1_MPORT_10_addr] <= ram_1_MPORT_10_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_11_en & ram_1_MPORT_11_mask) begin
      ram_1[ram_1_MPORT_11_addr] <= ram_1_MPORT_11_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_12_en & ram_1_MPORT_12_mask) begin
      ram_1[ram_1_MPORT_12_addr] <= ram_1_MPORT_12_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_13_en & ram_1_MPORT_13_mask) begin
      ram_1[ram_1_MPORT_13_addr] <= ram_1_MPORT_13_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_14_en & ram_1_MPORT_14_mask) begin
      ram_1[ram_1_MPORT_14_addr] <= ram_1_MPORT_14_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_15_en & ram_1_MPORT_15_mask) begin
      ram_1[ram_1_MPORT_15_addr] <= ram_1_MPORT_15_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_16_en & ram_1_MPORT_16_mask) begin
      ram_1[ram_1_MPORT_16_addr] <= ram_1_MPORT_16_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_17_en & ram_1_MPORT_17_mask) begin
      ram_1[ram_1_MPORT_17_addr] <= ram_1_MPORT_17_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_18_en & ram_1_MPORT_18_mask) begin
      ram_1[ram_1_MPORT_18_addr] <= ram_1_MPORT_18_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_19_en & ram_1_MPORT_19_mask) begin
      ram_1[ram_1_MPORT_19_addr] <= ram_1_MPORT_19_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_20_en & ram_1_MPORT_20_mask) begin
      ram_1[ram_1_MPORT_20_addr] <= ram_1_MPORT_20_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_21_en & ram_1_MPORT_21_mask) begin
      ram_1[ram_1_MPORT_21_addr] <= ram_1_MPORT_21_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_22_en & ram_1_MPORT_22_mask) begin
      ram_1[ram_1_MPORT_22_addr] <= ram_1_MPORT_22_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_23_en & ram_1_MPORT_23_mask) begin
      ram_1[ram_1_MPORT_23_addr] <= ram_1_MPORT_23_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_24_en & ram_1_MPORT_24_mask) begin
      ram_1[ram_1_MPORT_24_addr] <= ram_1_MPORT_24_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_25_en & ram_1_MPORT_25_mask) begin
      ram_1[ram_1_MPORT_25_addr] <= ram_1_MPORT_25_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_26_en & ram_1_MPORT_26_mask) begin
      ram_1[ram_1_MPORT_26_addr] <= ram_1_MPORT_26_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_27_en & ram_1_MPORT_27_mask) begin
      ram_1[ram_1_MPORT_27_addr] <= ram_1_MPORT_27_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_28_en & ram_1_MPORT_28_mask) begin
      ram_1[ram_1_MPORT_28_addr] <= ram_1_MPORT_28_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_29_en & ram_1_MPORT_29_mask) begin
      ram_1[ram_1_MPORT_29_addr] <= ram_1_MPORT_29_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_30_en & ram_1_MPORT_30_mask) begin
      ram_1[ram_1_MPORT_30_addr] <= ram_1_MPORT_30_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_31_en & ram_1_MPORT_31_mask) begin
      ram_1[ram_1_MPORT_31_addr] <= ram_1_MPORT_31_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_32_en & ram_1_MPORT_32_mask) begin
      ram_1[ram_1_MPORT_32_addr] <= ram_1_MPORT_32_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_33_en & ram_1_MPORT_33_mask) begin
      ram_1[ram_1_MPORT_33_addr] <= ram_1_MPORT_33_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_34_en & ram_1_MPORT_34_mask) begin
      ram_1[ram_1_MPORT_34_addr] <= ram_1_MPORT_34_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_35_en & ram_1_MPORT_35_mask) begin
      ram_1[ram_1_MPORT_35_addr] <= ram_1_MPORT_35_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_36_en & ram_1_MPORT_36_mask) begin
      ram_1[ram_1_MPORT_36_addr] <= ram_1_MPORT_36_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_37_en & ram_1_MPORT_37_mask) begin
      ram_1[ram_1_MPORT_37_addr] <= ram_1_MPORT_37_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_38_en & ram_1_MPORT_38_mask) begin
      ram_1[ram_1_MPORT_38_addr] <= ram_1_MPORT_38_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_39_en & ram_1_MPORT_39_mask) begin
      ram_1[ram_1_MPORT_39_addr] <= ram_1_MPORT_39_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_40_en & ram_1_MPORT_40_mask) begin
      ram_1[ram_1_MPORT_40_addr] <= ram_1_MPORT_40_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_41_en & ram_1_MPORT_41_mask) begin
      ram_1[ram_1_MPORT_41_addr] <= ram_1_MPORT_41_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_42_en & ram_1_MPORT_42_mask) begin
      ram_1[ram_1_MPORT_42_addr] <= ram_1_MPORT_42_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_43_en & ram_1_MPORT_43_mask) begin
      ram_1[ram_1_MPORT_43_addr] <= ram_1_MPORT_43_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_44_en & ram_1_MPORT_44_mask) begin
      ram_1[ram_1_MPORT_44_addr] <= ram_1_MPORT_44_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_45_en & ram_1_MPORT_45_mask) begin
      ram_1[ram_1_MPORT_45_addr] <= ram_1_MPORT_45_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_46_en & ram_1_MPORT_46_mask) begin
      ram_1[ram_1_MPORT_46_addr] <= ram_1_MPORT_46_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_47_en & ram_1_MPORT_47_mask) begin
      ram_1[ram_1_MPORT_47_addr] <= ram_1_MPORT_47_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_48_en & ram_1_MPORT_48_mask) begin
      ram_1[ram_1_MPORT_48_addr] <= ram_1_MPORT_48_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_49_en & ram_1_MPORT_49_mask) begin
      ram_1[ram_1_MPORT_49_addr] <= ram_1_MPORT_49_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_50_en & ram_1_MPORT_50_mask) begin
      ram_1[ram_1_MPORT_50_addr] <= ram_1_MPORT_50_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_51_en & ram_1_MPORT_51_mask) begin
      ram_1[ram_1_MPORT_51_addr] <= ram_1_MPORT_51_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_52_en & ram_1_MPORT_52_mask) begin
      ram_1[ram_1_MPORT_52_addr] <= ram_1_MPORT_52_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_53_en & ram_1_MPORT_53_mask) begin
      ram_1[ram_1_MPORT_53_addr] <= ram_1_MPORT_53_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_54_en & ram_1_MPORT_54_mask) begin
      ram_1[ram_1_MPORT_54_addr] <= ram_1_MPORT_54_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_55_en & ram_1_MPORT_55_mask) begin
      ram_1[ram_1_MPORT_55_addr] <= ram_1_MPORT_55_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_56_en & ram_1_MPORT_56_mask) begin
      ram_1[ram_1_MPORT_56_addr] <= ram_1_MPORT_56_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_57_en & ram_1_MPORT_57_mask) begin
      ram_1[ram_1_MPORT_57_addr] <= ram_1_MPORT_57_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_58_en & ram_1_MPORT_58_mask) begin
      ram_1[ram_1_MPORT_58_addr] <= ram_1_MPORT_58_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_59_en & ram_1_MPORT_59_mask) begin
      ram_1[ram_1_MPORT_59_addr] <= ram_1_MPORT_59_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_60_en & ram_1_MPORT_60_mask) begin
      ram_1[ram_1_MPORT_60_addr] <= ram_1_MPORT_60_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_61_en & ram_1_MPORT_61_mask) begin
      ram_1[ram_1_MPORT_61_addr] <= ram_1_MPORT_61_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_62_en & ram_1_MPORT_62_mask) begin
      ram_1[ram_1_MPORT_62_addr] <= ram_1_MPORT_62_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_63_en & ram_1_MPORT_63_mask) begin
      ram_1[ram_1_MPORT_63_addr] <= ram_1_MPORT_63_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_64_en & ram_1_MPORT_64_mask) begin
      ram_1[ram_1_MPORT_64_addr] <= ram_1_MPORT_64_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_65_en & ram_1_MPORT_65_mask) begin
      ram_1[ram_1_MPORT_65_addr] <= ram_1_MPORT_65_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_66_en & ram_1_MPORT_66_mask) begin
      ram_1[ram_1_MPORT_66_addr] <= ram_1_MPORT_66_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_67_en & ram_1_MPORT_67_mask) begin
      ram_1[ram_1_MPORT_67_addr] <= ram_1_MPORT_67_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_68_en & ram_1_MPORT_68_mask) begin
      ram_1[ram_1_MPORT_68_addr] <= ram_1_MPORT_68_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_69_en & ram_1_MPORT_69_mask) begin
      ram_1[ram_1_MPORT_69_addr] <= ram_1_MPORT_69_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_70_en & ram_1_MPORT_70_mask) begin
      ram_1[ram_1_MPORT_70_addr] <= ram_1_MPORT_70_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_71_en & ram_1_MPORT_71_mask) begin
      ram_1[ram_1_MPORT_71_addr] <= ram_1_MPORT_71_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_72_en & ram_1_MPORT_72_mask) begin
      ram_1[ram_1_MPORT_72_addr] <= ram_1_MPORT_72_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_73_en & ram_1_MPORT_73_mask) begin
      ram_1[ram_1_MPORT_73_addr] <= ram_1_MPORT_73_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_74_en & ram_1_MPORT_74_mask) begin
      ram_1[ram_1_MPORT_74_addr] <= ram_1_MPORT_74_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_75_en & ram_1_MPORT_75_mask) begin
      ram_1[ram_1_MPORT_75_addr] <= ram_1_MPORT_75_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_76_en & ram_1_MPORT_76_mask) begin
      ram_1[ram_1_MPORT_76_addr] <= ram_1_MPORT_76_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_77_en & ram_1_MPORT_77_mask) begin
      ram_1[ram_1_MPORT_77_addr] <= ram_1_MPORT_77_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_78_en & ram_1_MPORT_78_mask) begin
      ram_1[ram_1_MPORT_78_addr] <= ram_1_MPORT_78_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_79_en & ram_1_MPORT_79_mask) begin
      ram_1[ram_1_MPORT_79_addr] <= ram_1_MPORT_79_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_80_en & ram_1_MPORT_80_mask) begin
      ram_1[ram_1_MPORT_80_addr] <= ram_1_MPORT_80_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_81_en & ram_1_MPORT_81_mask) begin
      ram_1[ram_1_MPORT_81_addr] <= ram_1_MPORT_81_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_82_en & ram_1_MPORT_82_mask) begin
      ram_1[ram_1_MPORT_82_addr] <= ram_1_MPORT_82_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_83_en & ram_1_MPORT_83_mask) begin
      ram_1[ram_1_MPORT_83_addr] <= ram_1_MPORT_83_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_84_en & ram_1_MPORT_84_mask) begin
      ram_1[ram_1_MPORT_84_addr] <= ram_1_MPORT_84_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_85_en & ram_1_MPORT_85_mask) begin
      ram_1[ram_1_MPORT_85_addr] <= ram_1_MPORT_85_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_86_en & ram_1_MPORT_86_mask) begin
      ram_1[ram_1_MPORT_86_addr] <= ram_1_MPORT_86_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_87_en & ram_1_MPORT_87_mask) begin
      ram_1[ram_1_MPORT_87_addr] <= ram_1_MPORT_87_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_88_en & ram_1_MPORT_88_mask) begin
      ram_1[ram_1_MPORT_88_addr] <= ram_1_MPORT_88_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_89_en & ram_1_MPORT_89_mask) begin
      ram_1[ram_1_MPORT_89_addr] <= ram_1_MPORT_89_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_90_en & ram_1_MPORT_90_mask) begin
      ram_1[ram_1_MPORT_90_addr] <= ram_1_MPORT_90_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_91_en & ram_1_MPORT_91_mask) begin
      ram_1[ram_1_MPORT_91_addr] <= ram_1_MPORT_91_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_92_en & ram_1_MPORT_92_mask) begin
      ram_1[ram_1_MPORT_92_addr] <= ram_1_MPORT_92_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_93_en & ram_1_MPORT_93_mask) begin
      ram_1[ram_1_MPORT_93_addr] <= ram_1_MPORT_93_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_94_en & ram_1_MPORT_94_mask) begin
      ram_1[ram_1_MPORT_94_addr] <= ram_1_MPORT_94_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_95_en & ram_1_MPORT_95_mask) begin
      ram_1[ram_1_MPORT_95_addr] <= ram_1_MPORT_95_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_96_en & ram_1_MPORT_96_mask) begin
      ram_1[ram_1_MPORT_96_addr] <= ram_1_MPORT_96_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_97_en & ram_1_MPORT_97_mask) begin
      ram_1[ram_1_MPORT_97_addr] <= ram_1_MPORT_97_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_98_en & ram_1_MPORT_98_mask) begin
      ram_1[ram_1_MPORT_98_addr] <= ram_1_MPORT_98_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_99_en & ram_1_MPORT_99_mask) begin
      ram_1[ram_1_MPORT_99_addr] <= ram_1_MPORT_99_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_100_en & ram_1_MPORT_100_mask) begin
      ram_1[ram_1_MPORT_100_addr] <= ram_1_MPORT_100_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_101_en & ram_1_MPORT_101_mask) begin
      ram_1[ram_1_MPORT_101_addr] <= ram_1_MPORT_101_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_102_en & ram_1_MPORT_102_mask) begin
      ram_1[ram_1_MPORT_102_addr] <= ram_1_MPORT_102_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_103_en & ram_1_MPORT_103_mask) begin
      ram_1[ram_1_MPORT_103_addr] <= ram_1_MPORT_103_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_104_en & ram_1_MPORT_104_mask) begin
      ram_1[ram_1_MPORT_104_addr] <= ram_1_MPORT_104_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_105_en & ram_1_MPORT_105_mask) begin
      ram_1[ram_1_MPORT_105_addr] <= ram_1_MPORT_105_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_106_en & ram_1_MPORT_106_mask) begin
      ram_1[ram_1_MPORT_106_addr] <= ram_1_MPORT_106_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_107_en & ram_1_MPORT_107_mask) begin
      ram_1[ram_1_MPORT_107_addr] <= ram_1_MPORT_107_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_108_en & ram_1_MPORT_108_mask) begin
      ram_1[ram_1_MPORT_108_addr] <= ram_1_MPORT_108_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_109_en & ram_1_MPORT_109_mask) begin
      ram_1[ram_1_MPORT_109_addr] <= ram_1_MPORT_109_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_110_en & ram_1_MPORT_110_mask) begin
      ram_1[ram_1_MPORT_110_addr] <= ram_1_MPORT_110_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_111_en & ram_1_MPORT_111_mask) begin
      ram_1[ram_1_MPORT_111_addr] <= ram_1_MPORT_111_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_112_en & ram_1_MPORT_112_mask) begin
      ram_1[ram_1_MPORT_112_addr] <= ram_1_MPORT_112_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_113_en & ram_1_MPORT_113_mask) begin
      ram_1[ram_1_MPORT_113_addr] <= ram_1_MPORT_113_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_114_en & ram_1_MPORT_114_mask) begin
      ram_1[ram_1_MPORT_114_addr] <= ram_1_MPORT_114_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_115_en & ram_1_MPORT_115_mask) begin
      ram_1[ram_1_MPORT_115_addr] <= ram_1_MPORT_115_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_116_en & ram_1_MPORT_116_mask) begin
      ram_1[ram_1_MPORT_116_addr] <= ram_1_MPORT_116_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_117_en & ram_1_MPORT_117_mask) begin
      ram_1[ram_1_MPORT_117_addr] <= ram_1_MPORT_117_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_118_en & ram_1_MPORT_118_mask) begin
      ram_1[ram_1_MPORT_118_addr] <= ram_1_MPORT_118_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_119_en & ram_1_MPORT_119_mask) begin
      ram_1[ram_1_MPORT_119_addr] <= ram_1_MPORT_119_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_120_en & ram_1_MPORT_120_mask) begin
      ram_1[ram_1_MPORT_120_addr] <= ram_1_MPORT_120_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_121_en & ram_1_MPORT_121_mask) begin
      ram_1[ram_1_MPORT_121_addr] <= ram_1_MPORT_121_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_122_en & ram_1_MPORT_122_mask) begin
      ram_1[ram_1_MPORT_122_addr] <= ram_1_MPORT_122_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_123_en & ram_1_MPORT_123_mask) begin
      ram_1[ram_1_MPORT_123_addr] <= ram_1_MPORT_123_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_124_en & ram_1_MPORT_124_mask) begin
      ram_1[ram_1_MPORT_124_addr] <= ram_1_MPORT_124_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_125_en & ram_1_MPORT_125_mask) begin
      ram_1[ram_1_MPORT_125_addr] <= ram_1_MPORT_125_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_126_en & ram_1_MPORT_126_mask) begin
      ram_1[ram_1_MPORT_126_addr] <= ram_1_MPORT_126_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_127_en & ram_1_MPORT_127_mask) begin
      ram_1[ram_1_MPORT_127_addr] <= ram_1_MPORT_127_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_128_en & ram_1_MPORT_128_mask) begin
      ram_1[ram_1_MPORT_128_addr] <= ram_1_MPORT_128_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_129_en & ram_1_MPORT_129_mask) begin
      ram_1[ram_1_MPORT_129_addr] <= ram_1_MPORT_129_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_130_en & ram_1_MPORT_130_mask) begin
      ram_1[ram_1_MPORT_130_addr] <= ram_1_MPORT_130_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_131_en & ram_1_MPORT_131_mask) begin
      ram_1[ram_1_MPORT_131_addr] <= ram_1_MPORT_131_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_132_en & ram_1_MPORT_132_mask) begin
      ram_1[ram_1_MPORT_132_addr] <= ram_1_MPORT_132_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_133_en & ram_1_MPORT_133_mask) begin
      ram_1[ram_1_MPORT_133_addr] <= ram_1_MPORT_133_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_134_en & ram_1_MPORT_134_mask) begin
      ram_1[ram_1_MPORT_134_addr] <= ram_1_MPORT_134_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_135_en & ram_1_MPORT_135_mask) begin
      ram_1[ram_1_MPORT_135_addr] <= ram_1_MPORT_135_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_136_en & ram_1_MPORT_136_mask) begin
      ram_1[ram_1_MPORT_136_addr] <= ram_1_MPORT_136_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_137_en & ram_1_MPORT_137_mask) begin
      ram_1[ram_1_MPORT_137_addr] <= ram_1_MPORT_137_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_138_en & ram_1_MPORT_138_mask) begin
      ram_1[ram_1_MPORT_138_addr] <= ram_1_MPORT_138_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_139_en & ram_1_MPORT_139_mask) begin
      ram_1[ram_1_MPORT_139_addr] <= ram_1_MPORT_139_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_140_en & ram_1_MPORT_140_mask) begin
      ram_1[ram_1_MPORT_140_addr] <= ram_1_MPORT_140_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_141_en & ram_1_MPORT_141_mask) begin
      ram_1[ram_1_MPORT_141_addr] <= ram_1_MPORT_141_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_142_en & ram_1_MPORT_142_mask) begin
      ram_1[ram_1_MPORT_142_addr] <= ram_1_MPORT_142_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_143_en & ram_1_MPORT_143_mask) begin
      ram_1[ram_1_MPORT_143_addr] <= ram_1_MPORT_143_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_144_en & ram_1_MPORT_144_mask) begin
      ram_1[ram_1_MPORT_144_addr] <= ram_1_MPORT_144_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_145_en & ram_1_MPORT_145_mask) begin
      ram_1[ram_1_MPORT_145_addr] <= ram_1_MPORT_145_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_146_en & ram_1_MPORT_146_mask) begin
      ram_1[ram_1_MPORT_146_addr] <= ram_1_MPORT_146_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_147_en & ram_1_MPORT_147_mask) begin
      ram_1[ram_1_MPORT_147_addr] <= ram_1_MPORT_147_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_148_en & ram_1_MPORT_148_mask) begin
      ram_1[ram_1_MPORT_148_addr] <= ram_1_MPORT_148_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_149_en & ram_1_MPORT_149_mask) begin
      ram_1[ram_1_MPORT_149_addr] <= ram_1_MPORT_149_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_150_en & ram_1_MPORT_150_mask) begin
      ram_1[ram_1_MPORT_150_addr] <= ram_1_MPORT_150_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_151_en & ram_1_MPORT_151_mask) begin
      ram_1[ram_1_MPORT_151_addr] <= ram_1_MPORT_151_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_152_en & ram_1_MPORT_152_mask) begin
      ram_1[ram_1_MPORT_152_addr] <= ram_1_MPORT_152_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_153_en & ram_1_MPORT_153_mask) begin
      ram_1[ram_1_MPORT_153_addr] <= ram_1_MPORT_153_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_154_en & ram_1_MPORT_154_mask) begin
      ram_1[ram_1_MPORT_154_addr] <= ram_1_MPORT_154_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_155_en & ram_1_MPORT_155_mask) begin
      ram_1[ram_1_MPORT_155_addr] <= ram_1_MPORT_155_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_156_en & ram_1_MPORT_156_mask) begin
      ram_1[ram_1_MPORT_156_addr] <= ram_1_MPORT_156_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_157_en & ram_1_MPORT_157_mask) begin
      ram_1[ram_1_MPORT_157_addr] <= ram_1_MPORT_157_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_158_en & ram_1_MPORT_158_mask) begin
      ram_1[ram_1_MPORT_158_addr] <= ram_1_MPORT_158_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_159_en & ram_1_MPORT_159_mask) begin
      ram_1[ram_1_MPORT_159_addr] <= ram_1_MPORT_159_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_160_en & ram_1_MPORT_160_mask) begin
      ram_1[ram_1_MPORT_160_addr] <= ram_1_MPORT_160_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_161_en & ram_1_MPORT_161_mask) begin
      ram_1[ram_1_MPORT_161_addr] <= ram_1_MPORT_161_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_162_en & ram_1_MPORT_162_mask) begin
      ram_1[ram_1_MPORT_162_addr] <= ram_1_MPORT_162_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_163_en & ram_1_MPORT_163_mask) begin
      ram_1[ram_1_MPORT_163_addr] <= ram_1_MPORT_163_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_164_en & ram_1_MPORT_164_mask) begin
      ram_1[ram_1_MPORT_164_addr] <= ram_1_MPORT_164_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_165_en & ram_1_MPORT_165_mask) begin
      ram_1[ram_1_MPORT_165_addr] <= ram_1_MPORT_165_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_166_en & ram_1_MPORT_166_mask) begin
      ram_1[ram_1_MPORT_166_addr] <= ram_1_MPORT_166_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_167_en & ram_1_MPORT_167_mask) begin
      ram_1[ram_1_MPORT_167_addr] <= ram_1_MPORT_167_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_168_en & ram_1_MPORT_168_mask) begin
      ram_1[ram_1_MPORT_168_addr] <= ram_1_MPORT_168_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_169_en & ram_1_MPORT_169_mask) begin
      ram_1[ram_1_MPORT_169_addr] <= ram_1_MPORT_169_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_170_en & ram_1_MPORT_170_mask) begin
      ram_1[ram_1_MPORT_170_addr] <= ram_1_MPORT_170_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_171_en & ram_1_MPORT_171_mask) begin
      ram_1[ram_1_MPORT_171_addr] <= ram_1_MPORT_171_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_172_en & ram_1_MPORT_172_mask) begin
      ram_1[ram_1_MPORT_172_addr] <= ram_1_MPORT_172_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_173_en & ram_1_MPORT_173_mask) begin
      ram_1[ram_1_MPORT_173_addr] <= ram_1_MPORT_173_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_174_en & ram_1_MPORT_174_mask) begin
      ram_1[ram_1_MPORT_174_addr] <= ram_1_MPORT_174_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_175_en & ram_1_MPORT_175_mask) begin
      ram_1[ram_1_MPORT_175_addr] <= ram_1_MPORT_175_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_176_en & ram_1_MPORT_176_mask) begin
      ram_1[ram_1_MPORT_176_addr] <= ram_1_MPORT_176_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_177_en & ram_1_MPORT_177_mask) begin
      ram_1[ram_1_MPORT_177_addr] <= ram_1_MPORT_177_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_178_en & ram_1_MPORT_178_mask) begin
      ram_1[ram_1_MPORT_178_addr] <= ram_1_MPORT_178_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_179_en & ram_1_MPORT_179_mask) begin
      ram_1[ram_1_MPORT_179_addr] <= ram_1_MPORT_179_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_180_en & ram_1_MPORT_180_mask) begin
      ram_1[ram_1_MPORT_180_addr] <= ram_1_MPORT_180_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_181_en & ram_1_MPORT_181_mask) begin
      ram_1[ram_1_MPORT_181_addr] <= ram_1_MPORT_181_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_182_en & ram_1_MPORT_182_mask) begin
      ram_1[ram_1_MPORT_182_addr] <= ram_1_MPORT_182_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_183_en & ram_1_MPORT_183_mask) begin
      ram_1[ram_1_MPORT_183_addr] <= ram_1_MPORT_183_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_184_en & ram_1_MPORT_184_mask) begin
      ram_1[ram_1_MPORT_184_addr] <= ram_1_MPORT_184_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_185_en & ram_1_MPORT_185_mask) begin
      ram_1[ram_1_MPORT_185_addr] <= ram_1_MPORT_185_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_186_en & ram_1_MPORT_186_mask) begin
      ram_1[ram_1_MPORT_186_addr] <= ram_1_MPORT_186_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_187_en & ram_1_MPORT_187_mask) begin
      ram_1[ram_1_MPORT_187_addr] <= ram_1_MPORT_187_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_188_en & ram_1_MPORT_188_mask) begin
      ram_1[ram_1_MPORT_188_addr] <= ram_1_MPORT_188_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_189_en & ram_1_MPORT_189_mask) begin
      ram_1[ram_1_MPORT_189_addr] <= ram_1_MPORT_189_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_190_en & ram_1_MPORT_190_mask) begin
      ram_1[ram_1_MPORT_190_addr] <= ram_1_MPORT_190_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_191_en & ram_1_MPORT_191_mask) begin
      ram_1[ram_1_MPORT_191_addr] <= ram_1_MPORT_191_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_192_en & ram_1_MPORT_192_mask) begin
      ram_1[ram_1_MPORT_192_addr] <= ram_1_MPORT_192_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_193_en & ram_1_MPORT_193_mask) begin
      ram_1[ram_1_MPORT_193_addr] <= ram_1_MPORT_193_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_194_en & ram_1_MPORT_194_mask) begin
      ram_1[ram_1_MPORT_194_addr] <= ram_1_MPORT_194_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_195_en & ram_1_MPORT_195_mask) begin
      ram_1[ram_1_MPORT_195_addr] <= ram_1_MPORT_195_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_196_en & ram_1_MPORT_196_mask) begin
      ram_1[ram_1_MPORT_196_addr] <= ram_1_MPORT_196_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_197_en & ram_1_MPORT_197_mask) begin
      ram_1[ram_1_MPORT_197_addr] <= ram_1_MPORT_197_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_198_en & ram_1_MPORT_198_mask) begin
      ram_1[ram_1_MPORT_198_addr] <= ram_1_MPORT_198_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_199_en & ram_1_MPORT_199_mask) begin
      ram_1[ram_1_MPORT_199_addr] <= ram_1_MPORT_199_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_200_en & ram_1_MPORT_200_mask) begin
      ram_1[ram_1_MPORT_200_addr] <= ram_1_MPORT_200_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_201_en & ram_1_MPORT_201_mask) begin
      ram_1[ram_1_MPORT_201_addr] <= ram_1_MPORT_201_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_202_en & ram_1_MPORT_202_mask) begin
      ram_1[ram_1_MPORT_202_addr] <= ram_1_MPORT_202_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_203_en & ram_1_MPORT_203_mask) begin
      ram_1[ram_1_MPORT_203_addr] <= ram_1_MPORT_203_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_204_en & ram_1_MPORT_204_mask) begin
      ram_1[ram_1_MPORT_204_addr] <= ram_1_MPORT_204_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_205_en & ram_1_MPORT_205_mask) begin
      ram_1[ram_1_MPORT_205_addr] <= ram_1_MPORT_205_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_206_en & ram_1_MPORT_206_mask) begin
      ram_1[ram_1_MPORT_206_addr] <= ram_1_MPORT_206_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_207_en & ram_1_MPORT_207_mask) begin
      ram_1[ram_1_MPORT_207_addr] <= ram_1_MPORT_207_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_208_en & ram_1_MPORT_208_mask) begin
      ram_1[ram_1_MPORT_208_addr] <= ram_1_MPORT_208_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_209_en & ram_1_MPORT_209_mask) begin
      ram_1[ram_1_MPORT_209_addr] <= ram_1_MPORT_209_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_210_en & ram_1_MPORT_210_mask) begin
      ram_1[ram_1_MPORT_210_addr] <= ram_1_MPORT_210_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_211_en & ram_1_MPORT_211_mask) begin
      ram_1[ram_1_MPORT_211_addr] <= ram_1_MPORT_211_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_212_en & ram_1_MPORT_212_mask) begin
      ram_1[ram_1_MPORT_212_addr] <= ram_1_MPORT_212_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_213_en & ram_1_MPORT_213_mask) begin
      ram_1[ram_1_MPORT_213_addr] <= ram_1_MPORT_213_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_214_en & ram_1_MPORT_214_mask) begin
      ram_1[ram_1_MPORT_214_addr] <= ram_1_MPORT_214_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_215_en & ram_1_MPORT_215_mask) begin
      ram_1[ram_1_MPORT_215_addr] <= ram_1_MPORT_215_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_216_en & ram_1_MPORT_216_mask) begin
      ram_1[ram_1_MPORT_216_addr] <= ram_1_MPORT_216_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_217_en & ram_1_MPORT_217_mask) begin
      ram_1[ram_1_MPORT_217_addr] <= ram_1_MPORT_217_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_218_en & ram_1_MPORT_218_mask) begin
      ram_1[ram_1_MPORT_218_addr] <= ram_1_MPORT_218_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_219_en & ram_1_MPORT_219_mask) begin
      ram_1[ram_1_MPORT_219_addr] <= ram_1_MPORT_219_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_220_en & ram_1_MPORT_220_mask) begin
      ram_1[ram_1_MPORT_220_addr] <= ram_1_MPORT_220_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_221_en & ram_1_MPORT_221_mask) begin
      ram_1[ram_1_MPORT_221_addr] <= ram_1_MPORT_221_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_222_en & ram_1_MPORT_222_mask) begin
      ram_1[ram_1_MPORT_222_addr] <= ram_1_MPORT_222_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_223_en & ram_1_MPORT_223_mask) begin
      ram_1[ram_1_MPORT_223_addr] <= ram_1_MPORT_223_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_224_en & ram_1_MPORT_224_mask) begin
      ram_1[ram_1_MPORT_224_addr] <= ram_1_MPORT_224_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_225_en & ram_1_MPORT_225_mask) begin
      ram_1[ram_1_MPORT_225_addr] <= ram_1_MPORT_225_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_226_en & ram_1_MPORT_226_mask) begin
      ram_1[ram_1_MPORT_226_addr] <= ram_1_MPORT_226_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_227_en & ram_1_MPORT_227_mask) begin
      ram_1[ram_1_MPORT_227_addr] <= ram_1_MPORT_227_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_228_en & ram_1_MPORT_228_mask) begin
      ram_1[ram_1_MPORT_228_addr] <= ram_1_MPORT_228_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_229_en & ram_1_MPORT_229_mask) begin
      ram_1[ram_1_MPORT_229_addr] <= ram_1_MPORT_229_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_230_en & ram_1_MPORT_230_mask) begin
      ram_1[ram_1_MPORT_230_addr] <= ram_1_MPORT_230_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_231_en & ram_1_MPORT_231_mask) begin
      ram_1[ram_1_MPORT_231_addr] <= ram_1_MPORT_231_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_232_en & ram_1_MPORT_232_mask) begin
      ram_1[ram_1_MPORT_232_addr] <= ram_1_MPORT_232_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_233_en & ram_1_MPORT_233_mask) begin
      ram_1[ram_1_MPORT_233_addr] <= ram_1_MPORT_233_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_234_en & ram_1_MPORT_234_mask) begin
      ram_1[ram_1_MPORT_234_addr] <= ram_1_MPORT_234_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_235_en & ram_1_MPORT_235_mask) begin
      ram_1[ram_1_MPORT_235_addr] <= ram_1_MPORT_235_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_236_en & ram_1_MPORT_236_mask) begin
      ram_1[ram_1_MPORT_236_addr] <= ram_1_MPORT_236_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_237_en & ram_1_MPORT_237_mask) begin
      ram_1[ram_1_MPORT_237_addr] <= ram_1_MPORT_237_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_238_en & ram_1_MPORT_238_mask) begin
      ram_1[ram_1_MPORT_238_addr] <= ram_1_MPORT_238_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_239_en & ram_1_MPORT_239_mask) begin
      ram_1[ram_1_MPORT_239_addr] <= ram_1_MPORT_239_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_240_en & ram_1_MPORT_240_mask) begin
      ram_1[ram_1_MPORT_240_addr] <= ram_1_MPORT_240_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_241_en & ram_1_MPORT_241_mask) begin
      ram_1[ram_1_MPORT_241_addr] <= ram_1_MPORT_241_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_242_en & ram_1_MPORT_242_mask) begin
      ram_1[ram_1_MPORT_242_addr] <= ram_1_MPORT_242_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_243_en & ram_1_MPORT_243_mask) begin
      ram_1[ram_1_MPORT_243_addr] <= ram_1_MPORT_243_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_244_en & ram_1_MPORT_244_mask) begin
      ram_1[ram_1_MPORT_244_addr] <= ram_1_MPORT_244_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_245_en & ram_1_MPORT_245_mask) begin
      ram_1[ram_1_MPORT_245_addr] <= ram_1_MPORT_245_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_246_en & ram_1_MPORT_246_mask) begin
      ram_1[ram_1_MPORT_246_addr] <= ram_1_MPORT_246_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_247_en & ram_1_MPORT_247_mask) begin
      ram_1[ram_1_MPORT_247_addr] <= ram_1_MPORT_247_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_248_en & ram_1_MPORT_248_mask) begin
      ram_1[ram_1_MPORT_248_addr] <= ram_1_MPORT_248_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_249_en & ram_1_MPORT_249_mask) begin
      ram_1[ram_1_MPORT_249_addr] <= ram_1_MPORT_249_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_250_en & ram_1_MPORT_250_mask) begin
      ram_1[ram_1_MPORT_250_addr] <= ram_1_MPORT_250_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_251_en & ram_1_MPORT_251_mask) begin
      ram_1[ram_1_MPORT_251_addr] <= ram_1_MPORT_251_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_252_en & ram_1_MPORT_252_mask) begin
      ram_1[ram_1_MPORT_252_addr] <= ram_1_MPORT_252_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_253_en & ram_1_MPORT_253_mask) begin
      ram_1[ram_1_MPORT_253_addr] <= ram_1_MPORT_253_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_254_en & ram_1_MPORT_254_mask) begin
      ram_1[ram_1_MPORT_254_addr] <= ram_1_MPORT_254_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_255_en & ram_1_MPORT_255_mask) begin
      ram_1[ram_1_MPORT_255_addr] <= ram_1_MPORT_255_data; // @[SRAM.scala 36:26]
    end
    if (ram_1_MPORT_256_en & ram_1_MPORT_256_mask) begin
      ram_1[ram_1_MPORT_256_addr] <= ram_1_MPORT_256_data; // @[SRAM.scala 36:26]
    end
    if (io_rw) begin
      ram_1_io_rdata_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      ram_1_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    end
    if (io_rw ? 1'h0 : 1'h1) begin
      ram_1_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
    if (ram_2_MPORT_en & ram_2_MPORT_mask) begin
      ram_2[ram_2_MPORT_addr] <= ram_2_MPORT_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_1_en & ram_2_MPORT_1_mask) begin
      ram_2[ram_2_MPORT_1_addr] <= ram_2_MPORT_1_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_2_en & ram_2_MPORT_2_mask) begin
      ram_2[ram_2_MPORT_2_addr] <= ram_2_MPORT_2_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_3_en & ram_2_MPORT_3_mask) begin
      ram_2[ram_2_MPORT_3_addr] <= ram_2_MPORT_3_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_4_en & ram_2_MPORT_4_mask) begin
      ram_2[ram_2_MPORT_4_addr] <= ram_2_MPORT_4_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_5_en & ram_2_MPORT_5_mask) begin
      ram_2[ram_2_MPORT_5_addr] <= ram_2_MPORT_5_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_6_en & ram_2_MPORT_6_mask) begin
      ram_2[ram_2_MPORT_6_addr] <= ram_2_MPORT_6_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_7_en & ram_2_MPORT_7_mask) begin
      ram_2[ram_2_MPORT_7_addr] <= ram_2_MPORT_7_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_8_en & ram_2_MPORT_8_mask) begin
      ram_2[ram_2_MPORT_8_addr] <= ram_2_MPORT_8_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_9_en & ram_2_MPORT_9_mask) begin
      ram_2[ram_2_MPORT_9_addr] <= ram_2_MPORT_9_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_10_en & ram_2_MPORT_10_mask) begin
      ram_2[ram_2_MPORT_10_addr] <= ram_2_MPORT_10_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_11_en & ram_2_MPORT_11_mask) begin
      ram_2[ram_2_MPORT_11_addr] <= ram_2_MPORT_11_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_12_en & ram_2_MPORT_12_mask) begin
      ram_2[ram_2_MPORT_12_addr] <= ram_2_MPORT_12_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_13_en & ram_2_MPORT_13_mask) begin
      ram_2[ram_2_MPORT_13_addr] <= ram_2_MPORT_13_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_14_en & ram_2_MPORT_14_mask) begin
      ram_2[ram_2_MPORT_14_addr] <= ram_2_MPORT_14_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_15_en & ram_2_MPORT_15_mask) begin
      ram_2[ram_2_MPORT_15_addr] <= ram_2_MPORT_15_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_16_en & ram_2_MPORT_16_mask) begin
      ram_2[ram_2_MPORT_16_addr] <= ram_2_MPORT_16_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_17_en & ram_2_MPORT_17_mask) begin
      ram_2[ram_2_MPORT_17_addr] <= ram_2_MPORT_17_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_18_en & ram_2_MPORT_18_mask) begin
      ram_2[ram_2_MPORT_18_addr] <= ram_2_MPORT_18_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_19_en & ram_2_MPORT_19_mask) begin
      ram_2[ram_2_MPORT_19_addr] <= ram_2_MPORT_19_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_20_en & ram_2_MPORT_20_mask) begin
      ram_2[ram_2_MPORT_20_addr] <= ram_2_MPORT_20_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_21_en & ram_2_MPORT_21_mask) begin
      ram_2[ram_2_MPORT_21_addr] <= ram_2_MPORT_21_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_22_en & ram_2_MPORT_22_mask) begin
      ram_2[ram_2_MPORT_22_addr] <= ram_2_MPORT_22_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_23_en & ram_2_MPORT_23_mask) begin
      ram_2[ram_2_MPORT_23_addr] <= ram_2_MPORT_23_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_24_en & ram_2_MPORT_24_mask) begin
      ram_2[ram_2_MPORT_24_addr] <= ram_2_MPORT_24_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_25_en & ram_2_MPORT_25_mask) begin
      ram_2[ram_2_MPORT_25_addr] <= ram_2_MPORT_25_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_26_en & ram_2_MPORT_26_mask) begin
      ram_2[ram_2_MPORT_26_addr] <= ram_2_MPORT_26_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_27_en & ram_2_MPORT_27_mask) begin
      ram_2[ram_2_MPORT_27_addr] <= ram_2_MPORT_27_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_28_en & ram_2_MPORT_28_mask) begin
      ram_2[ram_2_MPORT_28_addr] <= ram_2_MPORT_28_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_29_en & ram_2_MPORT_29_mask) begin
      ram_2[ram_2_MPORT_29_addr] <= ram_2_MPORT_29_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_30_en & ram_2_MPORT_30_mask) begin
      ram_2[ram_2_MPORT_30_addr] <= ram_2_MPORT_30_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_31_en & ram_2_MPORT_31_mask) begin
      ram_2[ram_2_MPORT_31_addr] <= ram_2_MPORT_31_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_32_en & ram_2_MPORT_32_mask) begin
      ram_2[ram_2_MPORT_32_addr] <= ram_2_MPORT_32_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_33_en & ram_2_MPORT_33_mask) begin
      ram_2[ram_2_MPORT_33_addr] <= ram_2_MPORT_33_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_34_en & ram_2_MPORT_34_mask) begin
      ram_2[ram_2_MPORT_34_addr] <= ram_2_MPORT_34_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_35_en & ram_2_MPORT_35_mask) begin
      ram_2[ram_2_MPORT_35_addr] <= ram_2_MPORT_35_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_36_en & ram_2_MPORT_36_mask) begin
      ram_2[ram_2_MPORT_36_addr] <= ram_2_MPORT_36_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_37_en & ram_2_MPORT_37_mask) begin
      ram_2[ram_2_MPORT_37_addr] <= ram_2_MPORT_37_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_38_en & ram_2_MPORT_38_mask) begin
      ram_2[ram_2_MPORT_38_addr] <= ram_2_MPORT_38_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_39_en & ram_2_MPORT_39_mask) begin
      ram_2[ram_2_MPORT_39_addr] <= ram_2_MPORT_39_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_40_en & ram_2_MPORT_40_mask) begin
      ram_2[ram_2_MPORT_40_addr] <= ram_2_MPORT_40_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_41_en & ram_2_MPORT_41_mask) begin
      ram_2[ram_2_MPORT_41_addr] <= ram_2_MPORT_41_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_42_en & ram_2_MPORT_42_mask) begin
      ram_2[ram_2_MPORT_42_addr] <= ram_2_MPORT_42_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_43_en & ram_2_MPORT_43_mask) begin
      ram_2[ram_2_MPORT_43_addr] <= ram_2_MPORT_43_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_44_en & ram_2_MPORT_44_mask) begin
      ram_2[ram_2_MPORT_44_addr] <= ram_2_MPORT_44_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_45_en & ram_2_MPORT_45_mask) begin
      ram_2[ram_2_MPORT_45_addr] <= ram_2_MPORT_45_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_46_en & ram_2_MPORT_46_mask) begin
      ram_2[ram_2_MPORT_46_addr] <= ram_2_MPORT_46_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_47_en & ram_2_MPORT_47_mask) begin
      ram_2[ram_2_MPORT_47_addr] <= ram_2_MPORT_47_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_48_en & ram_2_MPORT_48_mask) begin
      ram_2[ram_2_MPORT_48_addr] <= ram_2_MPORT_48_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_49_en & ram_2_MPORT_49_mask) begin
      ram_2[ram_2_MPORT_49_addr] <= ram_2_MPORT_49_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_50_en & ram_2_MPORT_50_mask) begin
      ram_2[ram_2_MPORT_50_addr] <= ram_2_MPORT_50_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_51_en & ram_2_MPORT_51_mask) begin
      ram_2[ram_2_MPORT_51_addr] <= ram_2_MPORT_51_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_52_en & ram_2_MPORT_52_mask) begin
      ram_2[ram_2_MPORT_52_addr] <= ram_2_MPORT_52_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_53_en & ram_2_MPORT_53_mask) begin
      ram_2[ram_2_MPORT_53_addr] <= ram_2_MPORT_53_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_54_en & ram_2_MPORT_54_mask) begin
      ram_2[ram_2_MPORT_54_addr] <= ram_2_MPORT_54_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_55_en & ram_2_MPORT_55_mask) begin
      ram_2[ram_2_MPORT_55_addr] <= ram_2_MPORT_55_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_56_en & ram_2_MPORT_56_mask) begin
      ram_2[ram_2_MPORT_56_addr] <= ram_2_MPORT_56_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_57_en & ram_2_MPORT_57_mask) begin
      ram_2[ram_2_MPORT_57_addr] <= ram_2_MPORT_57_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_58_en & ram_2_MPORT_58_mask) begin
      ram_2[ram_2_MPORT_58_addr] <= ram_2_MPORT_58_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_59_en & ram_2_MPORT_59_mask) begin
      ram_2[ram_2_MPORT_59_addr] <= ram_2_MPORT_59_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_60_en & ram_2_MPORT_60_mask) begin
      ram_2[ram_2_MPORT_60_addr] <= ram_2_MPORT_60_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_61_en & ram_2_MPORT_61_mask) begin
      ram_2[ram_2_MPORT_61_addr] <= ram_2_MPORT_61_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_62_en & ram_2_MPORT_62_mask) begin
      ram_2[ram_2_MPORT_62_addr] <= ram_2_MPORT_62_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_63_en & ram_2_MPORT_63_mask) begin
      ram_2[ram_2_MPORT_63_addr] <= ram_2_MPORT_63_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_64_en & ram_2_MPORT_64_mask) begin
      ram_2[ram_2_MPORT_64_addr] <= ram_2_MPORT_64_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_65_en & ram_2_MPORT_65_mask) begin
      ram_2[ram_2_MPORT_65_addr] <= ram_2_MPORT_65_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_66_en & ram_2_MPORT_66_mask) begin
      ram_2[ram_2_MPORT_66_addr] <= ram_2_MPORT_66_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_67_en & ram_2_MPORT_67_mask) begin
      ram_2[ram_2_MPORT_67_addr] <= ram_2_MPORT_67_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_68_en & ram_2_MPORT_68_mask) begin
      ram_2[ram_2_MPORT_68_addr] <= ram_2_MPORT_68_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_69_en & ram_2_MPORT_69_mask) begin
      ram_2[ram_2_MPORT_69_addr] <= ram_2_MPORT_69_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_70_en & ram_2_MPORT_70_mask) begin
      ram_2[ram_2_MPORT_70_addr] <= ram_2_MPORT_70_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_71_en & ram_2_MPORT_71_mask) begin
      ram_2[ram_2_MPORT_71_addr] <= ram_2_MPORT_71_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_72_en & ram_2_MPORT_72_mask) begin
      ram_2[ram_2_MPORT_72_addr] <= ram_2_MPORT_72_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_73_en & ram_2_MPORT_73_mask) begin
      ram_2[ram_2_MPORT_73_addr] <= ram_2_MPORT_73_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_74_en & ram_2_MPORT_74_mask) begin
      ram_2[ram_2_MPORT_74_addr] <= ram_2_MPORT_74_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_75_en & ram_2_MPORT_75_mask) begin
      ram_2[ram_2_MPORT_75_addr] <= ram_2_MPORT_75_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_76_en & ram_2_MPORT_76_mask) begin
      ram_2[ram_2_MPORT_76_addr] <= ram_2_MPORT_76_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_77_en & ram_2_MPORT_77_mask) begin
      ram_2[ram_2_MPORT_77_addr] <= ram_2_MPORT_77_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_78_en & ram_2_MPORT_78_mask) begin
      ram_2[ram_2_MPORT_78_addr] <= ram_2_MPORT_78_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_79_en & ram_2_MPORT_79_mask) begin
      ram_2[ram_2_MPORT_79_addr] <= ram_2_MPORT_79_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_80_en & ram_2_MPORT_80_mask) begin
      ram_2[ram_2_MPORT_80_addr] <= ram_2_MPORT_80_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_81_en & ram_2_MPORT_81_mask) begin
      ram_2[ram_2_MPORT_81_addr] <= ram_2_MPORT_81_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_82_en & ram_2_MPORT_82_mask) begin
      ram_2[ram_2_MPORT_82_addr] <= ram_2_MPORT_82_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_83_en & ram_2_MPORT_83_mask) begin
      ram_2[ram_2_MPORT_83_addr] <= ram_2_MPORT_83_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_84_en & ram_2_MPORT_84_mask) begin
      ram_2[ram_2_MPORT_84_addr] <= ram_2_MPORT_84_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_85_en & ram_2_MPORT_85_mask) begin
      ram_2[ram_2_MPORT_85_addr] <= ram_2_MPORT_85_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_86_en & ram_2_MPORT_86_mask) begin
      ram_2[ram_2_MPORT_86_addr] <= ram_2_MPORT_86_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_87_en & ram_2_MPORT_87_mask) begin
      ram_2[ram_2_MPORT_87_addr] <= ram_2_MPORT_87_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_88_en & ram_2_MPORT_88_mask) begin
      ram_2[ram_2_MPORT_88_addr] <= ram_2_MPORT_88_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_89_en & ram_2_MPORT_89_mask) begin
      ram_2[ram_2_MPORT_89_addr] <= ram_2_MPORT_89_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_90_en & ram_2_MPORT_90_mask) begin
      ram_2[ram_2_MPORT_90_addr] <= ram_2_MPORT_90_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_91_en & ram_2_MPORT_91_mask) begin
      ram_2[ram_2_MPORT_91_addr] <= ram_2_MPORT_91_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_92_en & ram_2_MPORT_92_mask) begin
      ram_2[ram_2_MPORT_92_addr] <= ram_2_MPORT_92_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_93_en & ram_2_MPORT_93_mask) begin
      ram_2[ram_2_MPORT_93_addr] <= ram_2_MPORT_93_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_94_en & ram_2_MPORT_94_mask) begin
      ram_2[ram_2_MPORT_94_addr] <= ram_2_MPORT_94_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_95_en & ram_2_MPORT_95_mask) begin
      ram_2[ram_2_MPORT_95_addr] <= ram_2_MPORT_95_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_96_en & ram_2_MPORT_96_mask) begin
      ram_2[ram_2_MPORT_96_addr] <= ram_2_MPORT_96_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_97_en & ram_2_MPORT_97_mask) begin
      ram_2[ram_2_MPORT_97_addr] <= ram_2_MPORT_97_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_98_en & ram_2_MPORT_98_mask) begin
      ram_2[ram_2_MPORT_98_addr] <= ram_2_MPORT_98_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_99_en & ram_2_MPORT_99_mask) begin
      ram_2[ram_2_MPORT_99_addr] <= ram_2_MPORT_99_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_100_en & ram_2_MPORT_100_mask) begin
      ram_2[ram_2_MPORT_100_addr] <= ram_2_MPORT_100_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_101_en & ram_2_MPORT_101_mask) begin
      ram_2[ram_2_MPORT_101_addr] <= ram_2_MPORT_101_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_102_en & ram_2_MPORT_102_mask) begin
      ram_2[ram_2_MPORT_102_addr] <= ram_2_MPORT_102_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_103_en & ram_2_MPORT_103_mask) begin
      ram_2[ram_2_MPORT_103_addr] <= ram_2_MPORT_103_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_104_en & ram_2_MPORT_104_mask) begin
      ram_2[ram_2_MPORT_104_addr] <= ram_2_MPORT_104_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_105_en & ram_2_MPORT_105_mask) begin
      ram_2[ram_2_MPORT_105_addr] <= ram_2_MPORT_105_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_106_en & ram_2_MPORT_106_mask) begin
      ram_2[ram_2_MPORT_106_addr] <= ram_2_MPORT_106_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_107_en & ram_2_MPORT_107_mask) begin
      ram_2[ram_2_MPORT_107_addr] <= ram_2_MPORT_107_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_108_en & ram_2_MPORT_108_mask) begin
      ram_2[ram_2_MPORT_108_addr] <= ram_2_MPORT_108_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_109_en & ram_2_MPORT_109_mask) begin
      ram_2[ram_2_MPORT_109_addr] <= ram_2_MPORT_109_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_110_en & ram_2_MPORT_110_mask) begin
      ram_2[ram_2_MPORT_110_addr] <= ram_2_MPORT_110_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_111_en & ram_2_MPORT_111_mask) begin
      ram_2[ram_2_MPORT_111_addr] <= ram_2_MPORT_111_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_112_en & ram_2_MPORT_112_mask) begin
      ram_2[ram_2_MPORT_112_addr] <= ram_2_MPORT_112_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_113_en & ram_2_MPORT_113_mask) begin
      ram_2[ram_2_MPORT_113_addr] <= ram_2_MPORT_113_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_114_en & ram_2_MPORT_114_mask) begin
      ram_2[ram_2_MPORT_114_addr] <= ram_2_MPORT_114_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_115_en & ram_2_MPORT_115_mask) begin
      ram_2[ram_2_MPORT_115_addr] <= ram_2_MPORT_115_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_116_en & ram_2_MPORT_116_mask) begin
      ram_2[ram_2_MPORT_116_addr] <= ram_2_MPORT_116_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_117_en & ram_2_MPORT_117_mask) begin
      ram_2[ram_2_MPORT_117_addr] <= ram_2_MPORT_117_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_118_en & ram_2_MPORT_118_mask) begin
      ram_2[ram_2_MPORT_118_addr] <= ram_2_MPORT_118_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_119_en & ram_2_MPORT_119_mask) begin
      ram_2[ram_2_MPORT_119_addr] <= ram_2_MPORT_119_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_120_en & ram_2_MPORT_120_mask) begin
      ram_2[ram_2_MPORT_120_addr] <= ram_2_MPORT_120_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_121_en & ram_2_MPORT_121_mask) begin
      ram_2[ram_2_MPORT_121_addr] <= ram_2_MPORT_121_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_122_en & ram_2_MPORT_122_mask) begin
      ram_2[ram_2_MPORT_122_addr] <= ram_2_MPORT_122_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_123_en & ram_2_MPORT_123_mask) begin
      ram_2[ram_2_MPORT_123_addr] <= ram_2_MPORT_123_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_124_en & ram_2_MPORT_124_mask) begin
      ram_2[ram_2_MPORT_124_addr] <= ram_2_MPORT_124_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_125_en & ram_2_MPORT_125_mask) begin
      ram_2[ram_2_MPORT_125_addr] <= ram_2_MPORT_125_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_126_en & ram_2_MPORT_126_mask) begin
      ram_2[ram_2_MPORT_126_addr] <= ram_2_MPORT_126_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_127_en & ram_2_MPORT_127_mask) begin
      ram_2[ram_2_MPORT_127_addr] <= ram_2_MPORT_127_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_128_en & ram_2_MPORT_128_mask) begin
      ram_2[ram_2_MPORT_128_addr] <= ram_2_MPORT_128_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_129_en & ram_2_MPORT_129_mask) begin
      ram_2[ram_2_MPORT_129_addr] <= ram_2_MPORT_129_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_130_en & ram_2_MPORT_130_mask) begin
      ram_2[ram_2_MPORT_130_addr] <= ram_2_MPORT_130_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_131_en & ram_2_MPORT_131_mask) begin
      ram_2[ram_2_MPORT_131_addr] <= ram_2_MPORT_131_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_132_en & ram_2_MPORT_132_mask) begin
      ram_2[ram_2_MPORT_132_addr] <= ram_2_MPORT_132_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_133_en & ram_2_MPORT_133_mask) begin
      ram_2[ram_2_MPORT_133_addr] <= ram_2_MPORT_133_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_134_en & ram_2_MPORT_134_mask) begin
      ram_2[ram_2_MPORT_134_addr] <= ram_2_MPORT_134_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_135_en & ram_2_MPORT_135_mask) begin
      ram_2[ram_2_MPORT_135_addr] <= ram_2_MPORT_135_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_136_en & ram_2_MPORT_136_mask) begin
      ram_2[ram_2_MPORT_136_addr] <= ram_2_MPORT_136_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_137_en & ram_2_MPORT_137_mask) begin
      ram_2[ram_2_MPORT_137_addr] <= ram_2_MPORT_137_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_138_en & ram_2_MPORT_138_mask) begin
      ram_2[ram_2_MPORT_138_addr] <= ram_2_MPORT_138_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_139_en & ram_2_MPORT_139_mask) begin
      ram_2[ram_2_MPORT_139_addr] <= ram_2_MPORT_139_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_140_en & ram_2_MPORT_140_mask) begin
      ram_2[ram_2_MPORT_140_addr] <= ram_2_MPORT_140_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_141_en & ram_2_MPORT_141_mask) begin
      ram_2[ram_2_MPORT_141_addr] <= ram_2_MPORT_141_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_142_en & ram_2_MPORT_142_mask) begin
      ram_2[ram_2_MPORT_142_addr] <= ram_2_MPORT_142_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_143_en & ram_2_MPORT_143_mask) begin
      ram_2[ram_2_MPORT_143_addr] <= ram_2_MPORT_143_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_144_en & ram_2_MPORT_144_mask) begin
      ram_2[ram_2_MPORT_144_addr] <= ram_2_MPORT_144_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_145_en & ram_2_MPORT_145_mask) begin
      ram_2[ram_2_MPORT_145_addr] <= ram_2_MPORT_145_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_146_en & ram_2_MPORT_146_mask) begin
      ram_2[ram_2_MPORT_146_addr] <= ram_2_MPORT_146_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_147_en & ram_2_MPORT_147_mask) begin
      ram_2[ram_2_MPORT_147_addr] <= ram_2_MPORT_147_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_148_en & ram_2_MPORT_148_mask) begin
      ram_2[ram_2_MPORT_148_addr] <= ram_2_MPORT_148_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_149_en & ram_2_MPORT_149_mask) begin
      ram_2[ram_2_MPORT_149_addr] <= ram_2_MPORT_149_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_150_en & ram_2_MPORT_150_mask) begin
      ram_2[ram_2_MPORT_150_addr] <= ram_2_MPORT_150_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_151_en & ram_2_MPORT_151_mask) begin
      ram_2[ram_2_MPORT_151_addr] <= ram_2_MPORT_151_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_152_en & ram_2_MPORT_152_mask) begin
      ram_2[ram_2_MPORT_152_addr] <= ram_2_MPORT_152_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_153_en & ram_2_MPORT_153_mask) begin
      ram_2[ram_2_MPORT_153_addr] <= ram_2_MPORT_153_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_154_en & ram_2_MPORT_154_mask) begin
      ram_2[ram_2_MPORT_154_addr] <= ram_2_MPORT_154_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_155_en & ram_2_MPORT_155_mask) begin
      ram_2[ram_2_MPORT_155_addr] <= ram_2_MPORT_155_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_156_en & ram_2_MPORT_156_mask) begin
      ram_2[ram_2_MPORT_156_addr] <= ram_2_MPORT_156_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_157_en & ram_2_MPORT_157_mask) begin
      ram_2[ram_2_MPORT_157_addr] <= ram_2_MPORT_157_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_158_en & ram_2_MPORT_158_mask) begin
      ram_2[ram_2_MPORT_158_addr] <= ram_2_MPORT_158_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_159_en & ram_2_MPORT_159_mask) begin
      ram_2[ram_2_MPORT_159_addr] <= ram_2_MPORT_159_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_160_en & ram_2_MPORT_160_mask) begin
      ram_2[ram_2_MPORT_160_addr] <= ram_2_MPORT_160_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_161_en & ram_2_MPORT_161_mask) begin
      ram_2[ram_2_MPORT_161_addr] <= ram_2_MPORT_161_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_162_en & ram_2_MPORT_162_mask) begin
      ram_2[ram_2_MPORT_162_addr] <= ram_2_MPORT_162_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_163_en & ram_2_MPORT_163_mask) begin
      ram_2[ram_2_MPORT_163_addr] <= ram_2_MPORT_163_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_164_en & ram_2_MPORT_164_mask) begin
      ram_2[ram_2_MPORT_164_addr] <= ram_2_MPORT_164_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_165_en & ram_2_MPORT_165_mask) begin
      ram_2[ram_2_MPORT_165_addr] <= ram_2_MPORT_165_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_166_en & ram_2_MPORT_166_mask) begin
      ram_2[ram_2_MPORT_166_addr] <= ram_2_MPORT_166_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_167_en & ram_2_MPORT_167_mask) begin
      ram_2[ram_2_MPORT_167_addr] <= ram_2_MPORT_167_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_168_en & ram_2_MPORT_168_mask) begin
      ram_2[ram_2_MPORT_168_addr] <= ram_2_MPORT_168_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_169_en & ram_2_MPORT_169_mask) begin
      ram_2[ram_2_MPORT_169_addr] <= ram_2_MPORT_169_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_170_en & ram_2_MPORT_170_mask) begin
      ram_2[ram_2_MPORT_170_addr] <= ram_2_MPORT_170_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_171_en & ram_2_MPORT_171_mask) begin
      ram_2[ram_2_MPORT_171_addr] <= ram_2_MPORT_171_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_172_en & ram_2_MPORT_172_mask) begin
      ram_2[ram_2_MPORT_172_addr] <= ram_2_MPORT_172_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_173_en & ram_2_MPORT_173_mask) begin
      ram_2[ram_2_MPORT_173_addr] <= ram_2_MPORT_173_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_174_en & ram_2_MPORT_174_mask) begin
      ram_2[ram_2_MPORT_174_addr] <= ram_2_MPORT_174_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_175_en & ram_2_MPORT_175_mask) begin
      ram_2[ram_2_MPORT_175_addr] <= ram_2_MPORT_175_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_176_en & ram_2_MPORT_176_mask) begin
      ram_2[ram_2_MPORT_176_addr] <= ram_2_MPORT_176_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_177_en & ram_2_MPORT_177_mask) begin
      ram_2[ram_2_MPORT_177_addr] <= ram_2_MPORT_177_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_178_en & ram_2_MPORT_178_mask) begin
      ram_2[ram_2_MPORT_178_addr] <= ram_2_MPORT_178_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_179_en & ram_2_MPORT_179_mask) begin
      ram_2[ram_2_MPORT_179_addr] <= ram_2_MPORT_179_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_180_en & ram_2_MPORT_180_mask) begin
      ram_2[ram_2_MPORT_180_addr] <= ram_2_MPORT_180_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_181_en & ram_2_MPORT_181_mask) begin
      ram_2[ram_2_MPORT_181_addr] <= ram_2_MPORT_181_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_182_en & ram_2_MPORT_182_mask) begin
      ram_2[ram_2_MPORT_182_addr] <= ram_2_MPORT_182_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_183_en & ram_2_MPORT_183_mask) begin
      ram_2[ram_2_MPORT_183_addr] <= ram_2_MPORT_183_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_184_en & ram_2_MPORT_184_mask) begin
      ram_2[ram_2_MPORT_184_addr] <= ram_2_MPORT_184_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_185_en & ram_2_MPORT_185_mask) begin
      ram_2[ram_2_MPORT_185_addr] <= ram_2_MPORT_185_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_186_en & ram_2_MPORT_186_mask) begin
      ram_2[ram_2_MPORT_186_addr] <= ram_2_MPORT_186_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_187_en & ram_2_MPORT_187_mask) begin
      ram_2[ram_2_MPORT_187_addr] <= ram_2_MPORT_187_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_188_en & ram_2_MPORT_188_mask) begin
      ram_2[ram_2_MPORT_188_addr] <= ram_2_MPORT_188_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_189_en & ram_2_MPORT_189_mask) begin
      ram_2[ram_2_MPORT_189_addr] <= ram_2_MPORT_189_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_190_en & ram_2_MPORT_190_mask) begin
      ram_2[ram_2_MPORT_190_addr] <= ram_2_MPORT_190_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_191_en & ram_2_MPORT_191_mask) begin
      ram_2[ram_2_MPORT_191_addr] <= ram_2_MPORT_191_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_192_en & ram_2_MPORT_192_mask) begin
      ram_2[ram_2_MPORT_192_addr] <= ram_2_MPORT_192_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_193_en & ram_2_MPORT_193_mask) begin
      ram_2[ram_2_MPORT_193_addr] <= ram_2_MPORT_193_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_194_en & ram_2_MPORT_194_mask) begin
      ram_2[ram_2_MPORT_194_addr] <= ram_2_MPORT_194_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_195_en & ram_2_MPORT_195_mask) begin
      ram_2[ram_2_MPORT_195_addr] <= ram_2_MPORT_195_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_196_en & ram_2_MPORT_196_mask) begin
      ram_2[ram_2_MPORT_196_addr] <= ram_2_MPORT_196_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_197_en & ram_2_MPORT_197_mask) begin
      ram_2[ram_2_MPORT_197_addr] <= ram_2_MPORT_197_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_198_en & ram_2_MPORT_198_mask) begin
      ram_2[ram_2_MPORT_198_addr] <= ram_2_MPORT_198_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_199_en & ram_2_MPORT_199_mask) begin
      ram_2[ram_2_MPORT_199_addr] <= ram_2_MPORT_199_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_200_en & ram_2_MPORT_200_mask) begin
      ram_2[ram_2_MPORT_200_addr] <= ram_2_MPORT_200_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_201_en & ram_2_MPORT_201_mask) begin
      ram_2[ram_2_MPORT_201_addr] <= ram_2_MPORT_201_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_202_en & ram_2_MPORT_202_mask) begin
      ram_2[ram_2_MPORT_202_addr] <= ram_2_MPORT_202_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_203_en & ram_2_MPORT_203_mask) begin
      ram_2[ram_2_MPORT_203_addr] <= ram_2_MPORT_203_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_204_en & ram_2_MPORT_204_mask) begin
      ram_2[ram_2_MPORT_204_addr] <= ram_2_MPORT_204_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_205_en & ram_2_MPORT_205_mask) begin
      ram_2[ram_2_MPORT_205_addr] <= ram_2_MPORT_205_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_206_en & ram_2_MPORT_206_mask) begin
      ram_2[ram_2_MPORT_206_addr] <= ram_2_MPORT_206_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_207_en & ram_2_MPORT_207_mask) begin
      ram_2[ram_2_MPORT_207_addr] <= ram_2_MPORT_207_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_208_en & ram_2_MPORT_208_mask) begin
      ram_2[ram_2_MPORT_208_addr] <= ram_2_MPORT_208_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_209_en & ram_2_MPORT_209_mask) begin
      ram_2[ram_2_MPORT_209_addr] <= ram_2_MPORT_209_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_210_en & ram_2_MPORT_210_mask) begin
      ram_2[ram_2_MPORT_210_addr] <= ram_2_MPORT_210_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_211_en & ram_2_MPORT_211_mask) begin
      ram_2[ram_2_MPORT_211_addr] <= ram_2_MPORT_211_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_212_en & ram_2_MPORT_212_mask) begin
      ram_2[ram_2_MPORT_212_addr] <= ram_2_MPORT_212_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_213_en & ram_2_MPORT_213_mask) begin
      ram_2[ram_2_MPORT_213_addr] <= ram_2_MPORT_213_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_214_en & ram_2_MPORT_214_mask) begin
      ram_2[ram_2_MPORT_214_addr] <= ram_2_MPORT_214_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_215_en & ram_2_MPORT_215_mask) begin
      ram_2[ram_2_MPORT_215_addr] <= ram_2_MPORT_215_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_216_en & ram_2_MPORT_216_mask) begin
      ram_2[ram_2_MPORT_216_addr] <= ram_2_MPORT_216_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_217_en & ram_2_MPORT_217_mask) begin
      ram_2[ram_2_MPORT_217_addr] <= ram_2_MPORT_217_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_218_en & ram_2_MPORT_218_mask) begin
      ram_2[ram_2_MPORT_218_addr] <= ram_2_MPORT_218_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_219_en & ram_2_MPORT_219_mask) begin
      ram_2[ram_2_MPORT_219_addr] <= ram_2_MPORT_219_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_220_en & ram_2_MPORT_220_mask) begin
      ram_2[ram_2_MPORT_220_addr] <= ram_2_MPORT_220_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_221_en & ram_2_MPORT_221_mask) begin
      ram_2[ram_2_MPORT_221_addr] <= ram_2_MPORT_221_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_222_en & ram_2_MPORT_222_mask) begin
      ram_2[ram_2_MPORT_222_addr] <= ram_2_MPORT_222_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_223_en & ram_2_MPORT_223_mask) begin
      ram_2[ram_2_MPORT_223_addr] <= ram_2_MPORT_223_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_224_en & ram_2_MPORT_224_mask) begin
      ram_2[ram_2_MPORT_224_addr] <= ram_2_MPORT_224_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_225_en & ram_2_MPORT_225_mask) begin
      ram_2[ram_2_MPORT_225_addr] <= ram_2_MPORT_225_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_226_en & ram_2_MPORT_226_mask) begin
      ram_2[ram_2_MPORT_226_addr] <= ram_2_MPORT_226_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_227_en & ram_2_MPORT_227_mask) begin
      ram_2[ram_2_MPORT_227_addr] <= ram_2_MPORT_227_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_228_en & ram_2_MPORT_228_mask) begin
      ram_2[ram_2_MPORT_228_addr] <= ram_2_MPORT_228_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_229_en & ram_2_MPORT_229_mask) begin
      ram_2[ram_2_MPORT_229_addr] <= ram_2_MPORT_229_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_230_en & ram_2_MPORT_230_mask) begin
      ram_2[ram_2_MPORT_230_addr] <= ram_2_MPORT_230_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_231_en & ram_2_MPORT_231_mask) begin
      ram_2[ram_2_MPORT_231_addr] <= ram_2_MPORT_231_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_232_en & ram_2_MPORT_232_mask) begin
      ram_2[ram_2_MPORT_232_addr] <= ram_2_MPORT_232_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_233_en & ram_2_MPORT_233_mask) begin
      ram_2[ram_2_MPORT_233_addr] <= ram_2_MPORT_233_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_234_en & ram_2_MPORT_234_mask) begin
      ram_2[ram_2_MPORT_234_addr] <= ram_2_MPORT_234_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_235_en & ram_2_MPORT_235_mask) begin
      ram_2[ram_2_MPORT_235_addr] <= ram_2_MPORT_235_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_236_en & ram_2_MPORT_236_mask) begin
      ram_2[ram_2_MPORT_236_addr] <= ram_2_MPORT_236_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_237_en & ram_2_MPORT_237_mask) begin
      ram_2[ram_2_MPORT_237_addr] <= ram_2_MPORT_237_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_238_en & ram_2_MPORT_238_mask) begin
      ram_2[ram_2_MPORT_238_addr] <= ram_2_MPORT_238_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_239_en & ram_2_MPORT_239_mask) begin
      ram_2[ram_2_MPORT_239_addr] <= ram_2_MPORT_239_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_240_en & ram_2_MPORT_240_mask) begin
      ram_2[ram_2_MPORT_240_addr] <= ram_2_MPORT_240_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_241_en & ram_2_MPORT_241_mask) begin
      ram_2[ram_2_MPORT_241_addr] <= ram_2_MPORT_241_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_242_en & ram_2_MPORT_242_mask) begin
      ram_2[ram_2_MPORT_242_addr] <= ram_2_MPORT_242_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_243_en & ram_2_MPORT_243_mask) begin
      ram_2[ram_2_MPORT_243_addr] <= ram_2_MPORT_243_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_244_en & ram_2_MPORT_244_mask) begin
      ram_2[ram_2_MPORT_244_addr] <= ram_2_MPORT_244_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_245_en & ram_2_MPORT_245_mask) begin
      ram_2[ram_2_MPORT_245_addr] <= ram_2_MPORT_245_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_246_en & ram_2_MPORT_246_mask) begin
      ram_2[ram_2_MPORT_246_addr] <= ram_2_MPORT_246_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_247_en & ram_2_MPORT_247_mask) begin
      ram_2[ram_2_MPORT_247_addr] <= ram_2_MPORT_247_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_248_en & ram_2_MPORT_248_mask) begin
      ram_2[ram_2_MPORT_248_addr] <= ram_2_MPORT_248_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_249_en & ram_2_MPORT_249_mask) begin
      ram_2[ram_2_MPORT_249_addr] <= ram_2_MPORT_249_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_250_en & ram_2_MPORT_250_mask) begin
      ram_2[ram_2_MPORT_250_addr] <= ram_2_MPORT_250_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_251_en & ram_2_MPORT_251_mask) begin
      ram_2[ram_2_MPORT_251_addr] <= ram_2_MPORT_251_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_252_en & ram_2_MPORT_252_mask) begin
      ram_2[ram_2_MPORT_252_addr] <= ram_2_MPORT_252_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_253_en & ram_2_MPORT_253_mask) begin
      ram_2[ram_2_MPORT_253_addr] <= ram_2_MPORT_253_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_254_en & ram_2_MPORT_254_mask) begin
      ram_2[ram_2_MPORT_254_addr] <= ram_2_MPORT_254_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_255_en & ram_2_MPORT_255_mask) begin
      ram_2[ram_2_MPORT_255_addr] <= ram_2_MPORT_255_data; // @[SRAM.scala 36:26]
    end
    if (ram_2_MPORT_256_en & ram_2_MPORT_256_mask) begin
      ram_2[ram_2_MPORT_256_addr] <= ram_2_MPORT_256_data; // @[SRAM.scala 36:26]
    end
    if (io_rw) begin
      ram_2_io_rdata_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      ram_2_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    end
    if (io_rw ? 1'h0 : 1'h1) begin
      ram_2_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
    if (ram_3_MPORT_en & ram_3_MPORT_mask) begin
      ram_3[ram_3_MPORT_addr] <= ram_3_MPORT_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_1_en & ram_3_MPORT_1_mask) begin
      ram_3[ram_3_MPORT_1_addr] <= ram_3_MPORT_1_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_2_en & ram_3_MPORT_2_mask) begin
      ram_3[ram_3_MPORT_2_addr] <= ram_3_MPORT_2_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_3_en & ram_3_MPORT_3_mask) begin
      ram_3[ram_3_MPORT_3_addr] <= ram_3_MPORT_3_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_4_en & ram_3_MPORT_4_mask) begin
      ram_3[ram_3_MPORT_4_addr] <= ram_3_MPORT_4_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_5_en & ram_3_MPORT_5_mask) begin
      ram_3[ram_3_MPORT_5_addr] <= ram_3_MPORT_5_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_6_en & ram_3_MPORT_6_mask) begin
      ram_3[ram_3_MPORT_6_addr] <= ram_3_MPORT_6_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_7_en & ram_3_MPORT_7_mask) begin
      ram_3[ram_3_MPORT_7_addr] <= ram_3_MPORT_7_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_8_en & ram_3_MPORT_8_mask) begin
      ram_3[ram_3_MPORT_8_addr] <= ram_3_MPORT_8_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_9_en & ram_3_MPORT_9_mask) begin
      ram_3[ram_3_MPORT_9_addr] <= ram_3_MPORT_9_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_10_en & ram_3_MPORT_10_mask) begin
      ram_3[ram_3_MPORT_10_addr] <= ram_3_MPORT_10_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_11_en & ram_3_MPORT_11_mask) begin
      ram_3[ram_3_MPORT_11_addr] <= ram_3_MPORT_11_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_12_en & ram_3_MPORT_12_mask) begin
      ram_3[ram_3_MPORT_12_addr] <= ram_3_MPORT_12_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_13_en & ram_3_MPORT_13_mask) begin
      ram_3[ram_3_MPORT_13_addr] <= ram_3_MPORT_13_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_14_en & ram_3_MPORT_14_mask) begin
      ram_3[ram_3_MPORT_14_addr] <= ram_3_MPORT_14_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_15_en & ram_3_MPORT_15_mask) begin
      ram_3[ram_3_MPORT_15_addr] <= ram_3_MPORT_15_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_16_en & ram_3_MPORT_16_mask) begin
      ram_3[ram_3_MPORT_16_addr] <= ram_3_MPORT_16_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_17_en & ram_3_MPORT_17_mask) begin
      ram_3[ram_3_MPORT_17_addr] <= ram_3_MPORT_17_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_18_en & ram_3_MPORT_18_mask) begin
      ram_3[ram_3_MPORT_18_addr] <= ram_3_MPORT_18_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_19_en & ram_3_MPORT_19_mask) begin
      ram_3[ram_3_MPORT_19_addr] <= ram_3_MPORT_19_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_20_en & ram_3_MPORT_20_mask) begin
      ram_3[ram_3_MPORT_20_addr] <= ram_3_MPORT_20_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_21_en & ram_3_MPORT_21_mask) begin
      ram_3[ram_3_MPORT_21_addr] <= ram_3_MPORT_21_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_22_en & ram_3_MPORT_22_mask) begin
      ram_3[ram_3_MPORT_22_addr] <= ram_3_MPORT_22_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_23_en & ram_3_MPORT_23_mask) begin
      ram_3[ram_3_MPORT_23_addr] <= ram_3_MPORT_23_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_24_en & ram_3_MPORT_24_mask) begin
      ram_3[ram_3_MPORT_24_addr] <= ram_3_MPORT_24_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_25_en & ram_3_MPORT_25_mask) begin
      ram_3[ram_3_MPORT_25_addr] <= ram_3_MPORT_25_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_26_en & ram_3_MPORT_26_mask) begin
      ram_3[ram_3_MPORT_26_addr] <= ram_3_MPORT_26_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_27_en & ram_3_MPORT_27_mask) begin
      ram_3[ram_3_MPORT_27_addr] <= ram_3_MPORT_27_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_28_en & ram_3_MPORT_28_mask) begin
      ram_3[ram_3_MPORT_28_addr] <= ram_3_MPORT_28_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_29_en & ram_3_MPORT_29_mask) begin
      ram_3[ram_3_MPORT_29_addr] <= ram_3_MPORT_29_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_30_en & ram_3_MPORT_30_mask) begin
      ram_3[ram_3_MPORT_30_addr] <= ram_3_MPORT_30_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_31_en & ram_3_MPORT_31_mask) begin
      ram_3[ram_3_MPORT_31_addr] <= ram_3_MPORT_31_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_32_en & ram_3_MPORT_32_mask) begin
      ram_3[ram_3_MPORT_32_addr] <= ram_3_MPORT_32_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_33_en & ram_3_MPORT_33_mask) begin
      ram_3[ram_3_MPORT_33_addr] <= ram_3_MPORT_33_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_34_en & ram_3_MPORT_34_mask) begin
      ram_3[ram_3_MPORT_34_addr] <= ram_3_MPORT_34_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_35_en & ram_3_MPORT_35_mask) begin
      ram_3[ram_3_MPORT_35_addr] <= ram_3_MPORT_35_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_36_en & ram_3_MPORT_36_mask) begin
      ram_3[ram_3_MPORT_36_addr] <= ram_3_MPORT_36_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_37_en & ram_3_MPORT_37_mask) begin
      ram_3[ram_3_MPORT_37_addr] <= ram_3_MPORT_37_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_38_en & ram_3_MPORT_38_mask) begin
      ram_3[ram_3_MPORT_38_addr] <= ram_3_MPORT_38_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_39_en & ram_3_MPORT_39_mask) begin
      ram_3[ram_3_MPORT_39_addr] <= ram_3_MPORT_39_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_40_en & ram_3_MPORT_40_mask) begin
      ram_3[ram_3_MPORT_40_addr] <= ram_3_MPORT_40_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_41_en & ram_3_MPORT_41_mask) begin
      ram_3[ram_3_MPORT_41_addr] <= ram_3_MPORT_41_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_42_en & ram_3_MPORT_42_mask) begin
      ram_3[ram_3_MPORT_42_addr] <= ram_3_MPORT_42_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_43_en & ram_3_MPORT_43_mask) begin
      ram_3[ram_3_MPORT_43_addr] <= ram_3_MPORT_43_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_44_en & ram_3_MPORT_44_mask) begin
      ram_3[ram_3_MPORT_44_addr] <= ram_3_MPORT_44_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_45_en & ram_3_MPORT_45_mask) begin
      ram_3[ram_3_MPORT_45_addr] <= ram_3_MPORT_45_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_46_en & ram_3_MPORT_46_mask) begin
      ram_3[ram_3_MPORT_46_addr] <= ram_3_MPORT_46_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_47_en & ram_3_MPORT_47_mask) begin
      ram_3[ram_3_MPORT_47_addr] <= ram_3_MPORT_47_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_48_en & ram_3_MPORT_48_mask) begin
      ram_3[ram_3_MPORT_48_addr] <= ram_3_MPORT_48_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_49_en & ram_3_MPORT_49_mask) begin
      ram_3[ram_3_MPORT_49_addr] <= ram_3_MPORT_49_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_50_en & ram_3_MPORT_50_mask) begin
      ram_3[ram_3_MPORT_50_addr] <= ram_3_MPORT_50_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_51_en & ram_3_MPORT_51_mask) begin
      ram_3[ram_3_MPORT_51_addr] <= ram_3_MPORT_51_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_52_en & ram_3_MPORT_52_mask) begin
      ram_3[ram_3_MPORT_52_addr] <= ram_3_MPORT_52_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_53_en & ram_3_MPORT_53_mask) begin
      ram_3[ram_3_MPORT_53_addr] <= ram_3_MPORT_53_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_54_en & ram_3_MPORT_54_mask) begin
      ram_3[ram_3_MPORT_54_addr] <= ram_3_MPORT_54_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_55_en & ram_3_MPORT_55_mask) begin
      ram_3[ram_3_MPORT_55_addr] <= ram_3_MPORT_55_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_56_en & ram_3_MPORT_56_mask) begin
      ram_3[ram_3_MPORT_56_addr] <= ram_3_MPORT_56_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_57_en & ram_3_MPORT_57_mask) begin
      ram_3[ram_3_MPORT_57_addr] <= ram_3_MPORT_57_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_58_en & ram_3_MPORT_58_mask) begin
      ram_3[ram_3_MPORT_58_addr] <= ram_3_MPORT_58_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_59_en & ram_3_MPORT_59_mask) begin
      ram_3[ram_3_MPORT_59_addr] <= ram_3_MPORT_59_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_60_en & ram_3_MPORT_60_mask) begin
      ram_3[ram_3_MPORT_60_addr] <= ram_3_MPORT_60_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_61_en & ram_3_MPORT_61_mask) begin
      ram_3[ram_3_MPORT_61_addr] <= ram_3_MPORT_61_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_62_en & ram_3_MPORT_62_mask) begin
      ram_3[ram_3_MPORT_62_addr] <= ram_3_MPORT_62_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_63_en & ram_3_MPORT_63_mask) begin
      ram_3[ram_3_MPORT_63_addr] <= ram_3_MPORT_63_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_64_en & ram_3_MPORT_64_mask) begin
      ram_3[ram_3_MPORT_64_addr] <= ram_3_MPORT_64_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_65_en & ram_3_MPORT_65_mask) begin
      ram_3[ram_3_MPORT_65_addr] <= ram_3_MPORT_65_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_66_en & ram_3_MPORT_66_mask) begin
      ram_3[ram_3_MPORT_66_addr] <= ram_3_MPORT_66_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_67_en & ram_3_MPORT_67_mask) begin
      ram_3[ram_3_MPORT_67_addr] <= ram_3_MPORT_67_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_68_en & ram_3_MPORT_68_mask) begin
      ram_3[ram_3_MPORT_68_addr] <= ram_3_MPORT_68_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_69_en & ram_3_MPORT_69_mask) begin
      ram_3[ram_3_MPORT_69_addr] <= ram_3_MPORT_69_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_70_en & ram_3_MPORT_70_mask) begin
      ram_3[ram_3_MPORT_70_addr] <= ram_3_MPORT_70_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_71_en & ram_3_MPORT_71_mask) begin
      ram_3[ram_3_MPORT_71_addr] <= ram_3_MPORT_71_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_72_en & ram_3_MPORT_72_mask) begin
      ram_3[ram_3_MPORT_72_addr] <= ram_3_MPORT_72_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_73_en & ram_3_MPORT_73_mask) begin
      ram_3[ram_3_MPORT_73_addr] <= ram_3_MPORT_73_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_74_en & ram_3_MPORT_74_mask) begin
      ram_3[ram_3_MPORT_74_addr] <= ram_3_MPORT_74_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_75_en & ram_3_MPORT_75_mask) begin
      ram_3[ram_3_MPORT_75_addr] <= ram_3_MPORT_75_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_76_en & ram_3_MPORT_76_mask) begin
      ram_3[ram_3_MPORT_76_addr] <= ram_3_MPORT_76_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_77_en & ram_3_MPORT_77_mask) begin
      ram_3[ram_3_MPORT_77_addr] <= ram_3_MPORT_77_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_78_en & ram_3_MPORT_78_mask) begin
      ram_3[ram_3_MPORT_78_addr] <= ram_3_MPORT_78_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_79_en & ram_3_MPORT_79_mask) begin
      ram_3[ram_3_MPORT_79_addr] <= ram_3_MPORT_79_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_80_en & ram_3_MPORT_80_mask) begin
      ram_3[ram_3_MPORT_80_addr] <= ram_3_MPORT_80_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_81_en & ram_3_MPORT_81_mask) begin
      ram_3[ram_3_MPORT_81_addr] <= ram_3_MPORT_81_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_82_en & ram_3_MPORT_82_mask) begin
      ram_3[ram_3_MPORT_82_addr] <= ram_3_MPORT_82_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_83_en & ram_3_MPORT_83_mask) begin
      ram_3[ram_3_MPORT_83_addr] <= ram_3_MPORT_83_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_84_en & ram_3_MPORT_84_mask) begin
      ram_3[ram_3_MPORT_84_addr] <= ram_3_MPORT_84_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_85_en & ram_3_MPORT_85_mask) begin
      ram_3[ram_3_MPORT_85_addr] <= ram_3_MPORT_85_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_86_en & ram_3_MPORT_86_mask) begin
      ram_3[ram_3_MPORT_86_addr] <= ram_3_MPORT_86_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_87_en & ram_3_MPORT_87_mask) begin
      ram_3[ram_3_MPORT_87_addr] <= ram_3_MPORT_87_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_88_en & ram_3_MPORT_88_mask) begin
      ram_3[ram_3_MPORT_88_addr] <= ram_3_MPORT_88_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_89_en & ram_3_MPORT_89_mask) begin
      ram_3[ram_3_MPORT_89_addr] <= ram_3_MPORT_89_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_90_en & ram_3_MPORT_90_mask) begin
      ram_3[ram_3_MPORT_90_addr] <= ram_3_MPORT_90_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_91_en & ram_3_MPORT_91_mask) begin
      ram_3[ram_3_MPORT_91_addr] <= ram_3_MPORT_91_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_92_en & ram_3_MPORT_92_mask) begin
      ram_3[ram_3_MPORT_92_addr] <= ram_3_MPORT_92_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_93_en & ram_3_MPORT_93_mask) begin
      ram_3[ram_3_MPORT_93_addr] <= ram_3_MPORT_93_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_94_en & ram_3_MPORT_94_mask) begin
      ram_3[ram_3_MPORT_94_addr] <= ram_3_MPORT_94_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_95_en & ram_3_MPORT_95_mask) begin
      ram_3[ram_3_MPORT_95_addr] <= ram_3_MPORT_95_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_96_en & ram_3_MPORT_96_mask) begin
      ram_3[ram_3_MPORT_96_addr] <= ram_3_MPORT_96_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_97_en & ram_3_MPORT_97_mask) begin
      ram_3[ram_3_MPORT_97_addr] <= ram_3_MPORT_97_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_98_en & ram_3_MPORT_98_mask) begin
      ram_3[ram_3_MPORT_98_addr] <= ram_3_MPORT_98_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_99_en & ram_3_MPORT_99_mask) begin
      ram_3[ram_3_MPORT_99_addr] <= ram_3_MPORT_99_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_100_en & ram_3_MPORT_100_mask) begin
      ram_3[ram_3_MPORT_100_addr] <= ram_3_MPORT_100_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_101_en & ram_3_MPORT_101_mask) begin
      ram_3[ram_3_MPORT_101_addr] <= ram_3_MPORT_101_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_102_en & ram_3_MPORT_102_mask) begin
      ram_3[ram_3_MPORT_102_addr] <= ram_3_MPORT_102_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_103_en & ram_3_MPORT_103_mask) begin
      ram_3[ram_3_MPORT_103_addr] <= ram_3_MPORT_103_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_104_en & ram_3_MPORT_104_mask) begin
      ram_3[ram_3_MPORT_104_addr] <= ram_3_MPORT_104_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_105_en & ram_3_MPORT_105_mask) begin
      ram_3[ram_3_MPORT_105_addr] <= ram_3_MPORT_105_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_106_en & ram_3_MPORT_106_mask) begin
      ram_3[ram_3_MPORT_106_addr] <= ram_3_MPORT_106_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_107_en & ram_3_MPORT_107_mask) begin
      ram_3[ram_3_MPORT_107_addr] <= ram_3_MPORT_107_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_108_en & ram_3_MPORT_108_mask) begin
      ram_3[ram_3_MPORT_108_addr] <= ram_3_MPORT_108_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_109_en & ram_3_MPORT_109_mask) begin
      ram_3[ram_3_MPORT_109_addr] <= ram_3_MPORT_109_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_110_en & ram_3_MPORT_110_mask) begin
      ram_3[ram_3_MPORT_110_addr] <= ram_3_MPORT_110_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_111_en & ram_3_MPORT_111_mask) begin
      ram_3[ram_3_MPORT_111_addr] <= ram_3_MPORT_111_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_112_en & ram_3_MPORT_112_mask) begin
      ram_3[ram_3_MPORT_112_addr] <= ram_3_MPORT_112_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_113_en & ram_3_MPORT_113_mask) begin
      ram_3[ram_3_MPORT_113_addr] <= ram_3_MPORT_113_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_114_en & ram_3_MPORT_114_mask) begin
      ram_3[ram_3_MPORT_114_addr] <= ram_3_MPORT_114_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_115_en & ram_3_MPORT_115_mask) begin
      ram_3[ram_3_MPORT_115_addr] <= ram_3_MPORT_115_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_116_en & ram_3_MPORT_116_mask) begin
      ram_3[ram_3_MPORT_116_addr] <= ram_3_MPORT_116_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_117_en & ram_3_MPORT_117_mask) begin
      ram_3[ram_3_MPORT_117_addr] <= ram_3_MPORT_117_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_118_en & ram_3_MPORT_118_mask) begin
      ram_3[ram_3_MPORT_118_addr] <= ram_3_MPORT_118_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_119_en & ram_3_MPORT_119_mask) begin
      ram_3[ram_3_MPORT_119_addr] <= ram_3_MPORT_119_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_120_en & ram_3_MPORT_120_mask) begin
      ram_3[ram_3_MPORT_120_addr] <= ram_3_MPORT_120_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_121_en & ram_3_MPORT_121_mask) begin
      ram_3[ram_3_MPORT_121_addr] <= ram_3_MPORT_121_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_122_en & ram_3_MPORT_122_mask) begin
      ram_3[ram_3_MPORT_122_addr] <= ram_3_MPORT_122_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_123_en & ram_3_MPORT_123_mask) begin
      ram_3[ram_3_MPORT_123_addr] <= ram_3_MPORT_123_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_124_en & ram_3_MPORT_124_mask) begin
      ram_3[ram_3_MPORT_124_addr] <= ram_3_MPORT_124_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_125_en & ram_3_MPORT_125_mask) begin
      ram_3[ram_3_MPORT_125_addr] <= ram_3_MPORT_125_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_126_en & ram_3_MPORT_126_mask) begin
      ram_3[ram_3_MPORT_126_addr] <= ram_3_MPORT_126_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_127_en & ram_3_MPORT_127_mask) begin
      ram_3[ram_3_MPORT_127_addr] <= ram_3_MPORT_127_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_128_en & ram_3_MPORT_128_mask) begin
      ram_3[ram_3_MPORT_128_addr] <= ram_3_MPORT_128_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_129_en & ram_3_MPORT_129_mask) begin
      ram_3[ram_3_MPORT_129_addr] <= ram_3_MPORT_129_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_130_en & ram_3_MPORT_130_mask) begin
      ram_3[ram_3_MPORT_130_addr] <= ram_3_MPORT_130_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_131_en & ram_3_MPORT_131_mask) begin
      ram_3[ram_3_MPORT_131_addr] <= ram_3_MPORT_131_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_132_en & ram_3_MPORT_132_mask) begin
      ram_3[ram_3_MPORT_132_addr] <= ram_3_MPORT_132_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_133_en & ram_3_MPORT_133_mask) begin
      ram_3[ram_3_MPORT_133_addr] <= ram_3_MPORT_133_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_134_en & ram_3_MPORT_134_mask) begin
      ram_3[ram_3_MPORT_134_addr] <= ram_3_MPORT_134_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_135_en & ram_3_MPORT_135_mask) begin
      ram_3[ram_3_MPORT_135_addr] <= ram_3_MPORT_135_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_136_en & ram_3_MPORT_136_mask) begin
      ram_3[ram_3_MPORT_136_addr] <= ram_3_MPORT_136_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_137_en & ram_3_MPORT_137_mask) begin
      ram_3[ram_3_MPORT_137_addr] <= ram_3_MPORT_137_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_138_en & ram_3_MPORT_138_mask) begin
      ram_3[ram_3_MPORT_138_addr] <= ram_3_MPORT_138_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_139_en & ram_3_MPORT_139_mask) begin
      ram_3[ram_3_MPORT_139_addr] <= ram_3_MPORT_139_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_140_en & ram_3_MPORT_140_mask) begin
      ram_3[ram_3_MPORT_140_addr] <= ram_3_MPORT_140_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_141_en & ram_3_MPORT_141_mask) begin
      ram_3[ram_3_MPORT_141_addr] <= ram_3_MPORT_141_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_142_en & ram_3_MPORT_142_mask) begin
      ram_3[ram_3_MPORT_142_addr] <= ram_3_MPORT_142_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_143_en & ram_3_MPORT_143_mask) begin
      ram_3[ram_3_MPORT_143_addr] <= ram_3_MPORT_143_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_144_en & ram_3_MPORT_144_mask) begin
      ram_3[ram_3_MPORT_144_addr] <= ram_3_MPORT_144_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_145_en & ram_3_MPORT_145_mask) begin
      ram_3[ram_3_MPORT_145_addr] <= ram_3_MPORT_145_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_146_en & ram_3_MPORT_146_mask) begin
      ram_3[ram_3_MPORT_146_addr] <= ram_3_MPORT_146_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_147_en & ram_3_MPORT_147_mask) begin
      ram_3[ram_3_MPORT_147_addr] <= ram_3_MPORT_147_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_148_en & ram_3_MPORT_148_mask) begin
      ram_3[ram_3_MPORT_148_addr] <= ram_3_MPORT_148_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_149_en & ram_3_MPORT_149_mask) begin
      ram_3[ram_3_MPORT_149_addr] <= ram_3_MPORT_149_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_150_en & ram_3_MPORT_150_mask) begin
      ram_3[ram_3_MPORT_150_addr] <= ram_3_MPORT_150_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_151_en & ram_3_MPORT_151_mask) begin
      ram_3[ram_3_MPORT_151_addr] <= ram_3_MPORT_151_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_152_en & ram_3_MPORT_152_mask) begin
      ram_3[ram_3_MPORT_152_addr] <= ram_3_MPORT_152_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_153_en & ram_3_MPORT_153_mask) begin
      ram_3[ram_3_MPORT_153_addr] <= ram_3_MPORT_153_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_154_en & ram_3_MPORT_154_mask) begin
      ram_3[ram_3_MPORT_154_addr] <= ram_3_MPORT_154_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_155_en & ram_3_MPORT_155_mask) begin
      ram_3[ram_3_MPORT_155_addr] <= ram_3_MPORT_155_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_156_en & ram_3_MPORT_156_mask) begin
      ram_3[ram_3_MPORT_156_addr] <= ram_3_MPORT_156_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_157_en & ram_3_MPORT_157_mask) begin
      ram_3[ram_3_MPORT_157_addr] <= ram_3_MPORT_157_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_158_en & ram_3_MPORT_158_mask) begin
      ram_3[ram_3_MPORT_158_addr] <= ram_3_MPORT_158_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_159_en & ram_3_MPORT_159_mask) begin
      ram_3[ram_3_MPORT_159_addr] <= ram_3_MPORT_159_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_160_en & ram_3_MPORT_160_mask) begin
      ram_3[ram_3_MPORT_160_addr] <= ram_3_MPORT_160_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_161_en & ram_3_MPORT_161_mask) begin
      ram_3[ram_3_MPORT_161_addr] <= ram_3_MPORT_161_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_162_en & ram_3_MPORT_162_mask) begin
      ram_3[ram_3_MPORT_162_addr] <= ram_3_MPORT_162_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_163_en & ram_3_MPORT_163_mask) begin
      ram_3[ram_3_MPORT_163_addr] <= ram_3_MPORT_163_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_164_en & ram_3_MPORT_164_mask) begin
      ram_3[ram_3_MPORT_164_addr] <= ram_3_MPORT_164_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_165_en & ram_3_MPORT_165_mask) begin
      ram_3[ram_3_MPORT_165_addr] <= ram_3_MPORT_165_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_166_en & ram_3_MPORT_166_mask) begin
      ram_3[ram_3_MPORT_166_addr] <= ram_3_MPORT_166_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_167_en & ram_3_MPORT_167_mask) begin
      ram_3[ram_3_MPORT_167_addr] <= ram_3_MPORT_167_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_168_en & ram_3_MPORT_168_mask) begin
      ram_3[ram_3_MPORT_168_addr] <= ram_3_MPORT_168_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_169_en & ram_3_MPORT_169_mask) begin
      ram_3[ram_3_MPORT_169_addr] <= ram_3_MPORT_169_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_170_en & ram_3_MPORT_170_mask) begin
      ram_3[ram_3_MPORT_170_addr] <= ram_3_MPORT_170_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_171_en & ram_3_MPORT_171_mask) begin
      ram_3[ram_3_MPORT_171_addr] <= ram_3_MPORT_171_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_172_en & ram_3_MPORT_172_mask) begin
      ram_3[ram_3_MPORT_172_addr] <= ram_3_MPORT_172_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_173_en & ram_3_MPORT_173_mask) begin
      ram_3[ram_3_MPORT_173_addr] <= ram_3_MPORT_173_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_174_en & ram_3_MPORT_174_mask) begin
      ram_3[ram_3_MPORT_174_addr] <= ram_3_MPORT_174_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_175_en & ram_3_MPORT_175_mask) begin
      ram_3[ram_3_MPORT_175_addr] <= ram_3_MPORT_175_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_176_en & ram_3_MPORT_176_mask) begin
      ram_3[ram_3_MPORT_176_addr] <= ram_3_MPORT_176_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_177_en & ram_3_MPORT_177_mask) begin
      ram_3[ram_3_MPORT_177_addr] <= ram_3_MPORT_177_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_178_en & ram_3_MPORT_178_mask) begin
      ram_3[ram_3_MPORT_178_addr] <= ram_3_MPORT_178_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_179_en & ram_3_MPORT_179_mask) begin
      ram_3[ram_3_MPORT_179_addr] <= ram_3_MPORT_179_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_180_en & ram_3_MPORT_180_mask) begin
      ram_3[ram_3_MPORT_180_addr] <= ram_3_MPORT_180_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_181_en & ram_3_MPORT_181_mask) begin
      ram_3[ram_3_MPORT_181_addr] <= ram_3_MPORT_181_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_182_en & ram_3_MPORT_182_mask) begin
      ram_3[ram_3_MPORT_182_addr] <= ram_3_MPORT_182_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_183_en & ram_3_MPORT_183_mask) begin
      ram_3[ram_3_MPORT_183_addr] <= ram_3_MPORT_183_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_184_en & ram_3_MPORT_184_mask) begin
      ram_3[ram_3_MPORT_184_addr] <= ram_3_MPORT_184_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_185_en & ram_3_MPORT_185_mask) begin
      ram_3[ram_3_MPORT_185_addr] <= ram_3_MPORT_185_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_186_en & ram_3_MPORT_186_mask) begin
      ram_3[ram_3_MPORT_186_addr] <= ram_3_MPORT_186_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_187_en & ram_3_MPORT_187_mask) begin
      ram_3[ram_3_MPORT_187_addr] <= ram_3_MPORT_187_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_188_en & ram_3_MPORT_188_mask) begin
      ram_3[ram_3_MPORT_188_addr] <= ram_3_MPORT_188_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_189_en & ram_3_MPORT_189_mask) begin
      ram_3[ram_3_MPORT_189_addr] <= ram_3_MPORT_189_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_190_en & ram_3_MPORT_190_mask) begin
      ram_3[ram_3_MPORT_190_addr] <= ram_3_MPORT_190_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_191_en & ram_3_MPORT_191_mask) begin
      ram_3[ram_3_MPORT_191_addr] <= ram_3_MPORT_191_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_192_en & ram_3_MPORT_192_mask) begin
      ram_3[ram_3_MPORT_192_addr] <= ram_3_MPORT_192_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_193_en & ram_3_MPORT_193_mask) begin
      ram_3[ram_3_MPORT_193_addr] <= ram_3_MPORT_193_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_194_en & ram_3_MPORT_194_mask) begin
      ram_3[ram_3_MPORT_194_addr] <= ram_3_MPORT_194_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_195_en & ram_3_MPORT_195_mask) begin
      ram_3[ram_3_MPORT_195_addr] <= ram_3_MPORT_195_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_196_en & ram_3_MPORT_196_mask) begin
      ram_3[ram_3_MPORT_196_addr] <= ram_3_MPORT_196_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_197_en & ram_3_MPORT_197_mask) begin
      ram_3[ram_3_MPORT_197_addr] <= ram_3_MPORT_197_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_198_en & ram_3_MPORT_198_mask) begin
      ram_3[ram_3_MPORT_198_addr] <= ram_3_MPORT_198_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_199_en & ram_3_MPORT_199_mask) begin
      ram_3[ram_3_MPORT_199_addr] <= ram_3_MPORT_199_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_200_en & ram_3_MPORT_200_mask) begin
      ram_3[ram_3_MPORT_200_addr] <= ram_3_MPORT_200_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_201_en & ram_3_MPORT_201_mask) begin
      ram_3[ram_3_MPORT_201_addr] <= ram_3_MPORT_201_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_202_en & ram_3_MPORT_202_mask) begin
      ram_3[ram_3_MPORT_202_addr] <= ram_3_MPORT_202_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_203_en & ram_3_MPORT_203_mask) begin
      ram_3[ram_3_MPORT_203_addr] <= ram_3_MPORT_203_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_204_en & ram_3_MPORT_204_mask) begin
      ram_3[ram_3_MPORT_204_addr] <= ram_3_MPORT_204_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_205_en & ram_3_MPORT_205_mask) begin
      ram_3[ram_3_MPORT_205_addr] <= ram_3_MPORT_205_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_206_en & ram_3_MPORT_206_mask) begin
      ram_3[ram_3_MPORT_206_addr] <= ram_3_MPORT_206_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_207_en & ram_3_MPORT_207_mask) begin
      ram_3[ram_3_MPORT_207_addr] <= ram_3_MPORT_207_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_208_en & ram_3_MPORT_208_mask) begin
      ram_3[ram_3_MPORT_208_addr] <= ram_3_MPORT_208_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_209_en & ram_3_MPORT_209_mask) begin
      ram_3[ram_3_MPORT_209_addr] <= ram_3_MPORT_209_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_210_en & ram_3_MPORT_210_mask) begin
      ram_3[ram_3_MPORT_210_addr] <= ram_3_MPORT_210_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_211_en & ram_3_MPORT_211_mask) begin
      ram_3[ram_3_MPORT_211_addr] <= ram_3_MPORT_211_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_212_en & ram_3_MPORT_212_mask) begin
      ram_3[ram_3_MPORT_212_addr] <= ram_3_MPORT_212_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_213_en & ram_3_MPORT_213_mask) begin
      ram_3[ram_3_MPORT_213_addr] <= ram_3_MPORT_213_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_214_en & ram_3_MPORT_214_mask) begin
      ram_3[ram_3_MPORT_214_addr] <= ram_3_MPORT_214_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_215_en & ram_3_MPORT_215_mask) begin
      ram_3[ram_3_MPORT_215_addr] <= ram_3_MPORT_215_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_216_en & ram_3_MPORT_216_mask) begin
      ram_3[ram_3_MPORT_216_addr] <= ram_3_MPORT_216_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_217_en & ram_3_MPORT_217_mask) begin
      ram_3[ram_3_MPORT_217_addr] <= ram_3_MPORT_217_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_218_en & ram_3_MPORT_218_mask) begin
      ram_3[ram_3_MPORT_218_addr] <= ram_3_MPORT_218_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_219_en & ram_3_MPORT_219_mask) begin
      ram_3[ram_3_MPORT_219_addr] <= ram_3_MPORT_219_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_220_en & ram_3_MPORT_220_mask) begin
      ram_3[ram_3_MPORT_220_addr] <= ram_3_MPORT_220_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_221_en & ram_3_MPORT_221_mask) begin
      ram_3[ram_3_MPORT_221_addr] <= ram_3_MPORT_221_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_222_en & ram_3_MPORT_222_mask) begin
      ram_3[ram_3_MPORT_222_addr] <= ram_3_MPORT_222_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_223_en & ram_3_MPORT_223_mask) begin
      ram_3[ram_3_MPORT_223_addr] <= ram_3_MPORT_223_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_224_en & ram_3_MPORT_224_mask) begin
      ram_3[ram_3_MPORT_224_addr] <= ram_3_MPORT_224_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_225_en & ram_3_MPORT_225_mask) begin
      ram_3[ram_3_MPORT_225_addr] <= ram_3_MPORT_225_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_226_en & ram_3_MPORT_226_mask) begin
      ram_3[ram_3_MPORT_226_addr] <= ram_3_MPORT_226_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_227_en & ram_3_MPORT_227_mask) begin
      ram_3[ram_3_MPORT_227_addr] <= ram_3_MPORT_227_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_228_en & ram_3_MPORT_228_mask) begin
      ram_3[ram_3_MPORT_228_addr] <= ram_3_MPORT_228_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_229_en & ram_3_MPORT_229_mask) begin
      ram_3[ram_3_MPORT_229_addr] <= ram_3_MPORT_229_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_230_en & ram_3_MPORT_230_mask) begin
      ram_3[ram_3_MPORT_230_addr] <= ram_3_MPORT_230_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_231_en & ram_3_MPORT_231_mask) begin
      ram_3[ram_3_MPORT_231_addr] <= ram_3_MPORT_231_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_232_en & ram_3_MPORT_232_mask) begin
      ram_3[ram_3_MPORT_232_addr] <= ram_3_MPORT_232_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_233_en & ram_3_MPORT_233_mask) begin
      ram_3[ram_3_MPORT_233_addr] <= ram_3_MPORT_233_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_234_en & ram_3_MPORT_234_mask) begin
      ram_3[ram_3_MPORT_234_addr] <= ram_3_MPORT_234_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_235_en & ram_3_MPORT_235_mask) begin
      ram_3[ram_3_MPORT_235_addr] <= ram_3_MPORT_235_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_236_en & ram_3_MPORT_236_mask) begin
      ram_3[ram_3_MPORT_236_addr] <= ram_3_MPORT_236_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_237_en & ram_3_MPORT_237_mask) begin
      ram_3[ram_3_MPORT_237_addr] <= ram_3_MPORT_237_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_238_en & ram_3_MPORT_238_mask) begin
      ram_3[ram_3_MPORT_238_addr] <= ram_3_MPORT_238_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_239_en & ram_3_MPORT_239_mask) begin
      ram_3[ram_3_MPORT_239_addr] <= ram_3_MPORT_239_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_240_en & ram_3_MPORT_240_mask) begin
      ram_3[ram_3_MPORT_240_addr] <= ram_3_MPORT_240_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_241_en & ram_3_MPORT_241_mask) begin
      ram_3[ram_3_MPORT_241_addr] <= ram_3_MPORT_241_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_242_en & ram_3_MPORT_242_mask) begin
      ram_3[ram_3_MPORT_242_addr] <= ram_3_MPORT_242_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_243_en & ram_3_MPORT_243_mask) begin
      ram_3[ram_3_MPORT_243_addr] <= ram_3_MPORT_243_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_244_en & ram_3_MPORT_244_mask) begin
      ram_3[ram_3_MPORT_244_addr] <= ram_3_MPORT_244_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_245_en & ram_3_MPORT_245_mask) begin
      ram_3[ram_3_MPORT_245_addr] <= ram_3_MPORT_245_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_246_en & ram_3_MPORT_246_mask) begin
      ram_3[ram_3_MPORT_246_addr] <= ram_3_MPORT_246_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_247_en & ram_3_MPORT_247_mask) begin
      ram_3[ram_3_MPORT_247_addr] <= ram_3_MPORT_247_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_248_en & ram_3_MPORT_248_mask) begin
      ram_3[ram_3_MPORT_248_addr] <= ram_3_MPORT_248_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_249_en & ram_3_MPORT_249_mask) begin
      ram_3[ram_3_MPORT_249_addr] <= ram_3_MPORT_249_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_250_en & ram_3_MPORT_250_mask) begin
      ram_3[ram_3_MPORT_250_addr] <= ram_3_MPORT_250_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_251_en & ram_3_MPORT_251_mask) begin
      ram_3[ram_3_MPORT_251_addr] <= ram_3_MPORT_251_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_252_en & ram_3_MPORT_252_mask) begin
      ram_3[ram_3_MPORT_252_addr] <= ram_3_MPORT_252_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_253_en & ram_3_MPORT_253_mask) begin
      ram_3[ram_3_MPORT_253_addr] <= ram_3_MPORT_253_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_254_en & ram_3_MPORT_254_mask) begin
      ram_3[ram_3_MPORT_254_addr] <= ram_3_MPORT_254_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_255_en & ram_3_MPORT_255_mask) begin
      ram_3[ram_3_MPORT_255_addr] <= ram_3_MPORT_255_data; // @[SRAM.scala 36:26]
    end
    if (ram_3_MPORT_256_en & ram_3_MPORT_256_mask) begin
      ram_3[ram_3_MPORT_256_addr] <= ram_3_MPORT_256_data; // @[SRAM.scala 36:26]
    end
    if (io_rw) begin
      ram_3_io_rdata_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      ram_3_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    end
    if (io_rw ? 1'h0 : 1'h1) begin
      ram_3_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram_0[initvar] = _RAND_0[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram_1[initvar] = _RAND_3[1:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram_2[initvar] = _RAND_6[1:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram_3[initvar] = _RAND_9[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_0_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_0_io_rdata_MPORT_addr_pipe_0 = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  ram_1_io_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ram_1_io_rdata_MPORT_addr_pipe_0 = _RAND_5[7:0];
  _RAND_7 = {1{`RANDOM}};
  ram_2_io_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ram_2_io_rdata_MPORT_addr_pipe_0 = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  ram_3_io_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ram_3_io_rdata_MPORT_addr_pipe_0 = _RAND_11[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
