module BankRAM_2P(
  input         clock,
  input         reset,
  input  [6:0]  io_r_addr,
  output [31:0] io_r_data,
  input         io_w_en,
  input  [6:0]  io_w_addr,
  input  [31:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:127]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [6:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 32'h0;
  assign mem_MPORT_addr = 7'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 32'h0;
  assign mem_MPORT_1_addr = 7'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 32'h0;
  assign mem_MPORT_2_addr = 7'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 32'h0;
  assign mem_MPORT_3_addr = 7'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 32'h0;
  assign mem_MPORT_4_addr = 7'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 32'h0;
  assign mem_MPORT_5_addr = 7'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 32'h0;
  assign mem_MPORT_6_addr = 7'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 32'h0;
  assign mem_MPORT_7_addr = 7'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 32'h0;
  assign mem_MPORT_8_addr = 7'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 32'h0;
  assign mem_MPORT_9_addr = 7'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 32'h0;
  assign mem_MPORT_10_addr = 7'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 32'h0;
  assign mem_MPORT_11_addr = 7'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 32'h0;
  assign mem_MPORT_12_addr = 7'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 32'h0;
  assign mem_MPORT_13_addr = 7'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 32'h0;
  assign mem_MPORT_14_addr = 7'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 32'h0;
  assign mem_MPORT_15_addr = 7'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 32'h0;
  assign mem_MPORT_16_addr = 7'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 32'h0;
  assign mem_MPORT_17_addr = 7'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 32'h0;
  assign mem_MPORT_18_addr = 7'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 32'h0;
  assign mem_MPORT_19_addr = 7'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 32'h0;
  assign mem_MPORT_20_addr = 7'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 32'h0;
  assign mem_MPORT_21_addr = 7'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 32'h0;
  assign mem_MPORT_22_addr = 7'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 32'h0;
  assign mem_MPORT_23_addr = 7'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 32'h0;
  assign mem_MPORT_24_addr = 7'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 32'h0;
  assign mem_MPORT_25_addr = 7'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 32'h0;
  assign mem_MPORT_26_addr = 7'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 32'h0;
  assign mem_MPORT_27_addr = 7'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 32'h0;
  assign mem_MPORT_28_addr = 7'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 32'h0;
  assign mem_MPORT_29_addr = 7'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 32'h0;
  assign mem_MPORT_30_addr = 7'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 32'h0;
  assign mem_MPORT_31_addr = 7'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 32'h0;
  assign mem_MPORT_32_addr = 7'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 32'h0;
  assign mem_MPORT_33_addr = 7'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 32'h0;
  assign mem_MPORT_34_addr = 7'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 32'h0;
  assign mem_MPORT_35_addr = 7'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 32'h0;
  assign mem_MPORT_36_addr = 7'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 32'h0;
  assign mem_MPORT_37_addr = 7'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 32'h0;
  assign mem_MPORT_38_addr = 7'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 32'h0;
  assign mem_MPORT_39_addr = 7'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 32'h0;
  assign mem_MPORT_40_addr = 7'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 32'h0;
  assign mem_MPORT_41_addr = 7'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 32'h0;
  assign mem_MPORT_42_addr = 7'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 32'h0;
  assign mem_MPORT_43_addr = 7'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 32'h0;
  assign mem_MPORT_44_addr = 7'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 32'h0;
  assign mem_MPORT_45_addr = 7'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 32'h0;
  assign mem_MPORT_46_addr = 7'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 32'h0;
  assign mem_MPORT_47_addr = 7'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 32'h0;
  assign mem_MPORT_48_addr = 7'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 32'h0;
  assign mem_MPORT_49_addr = 7'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 32'h0;
  assign mem_MPORT_50_addr = 7'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 32'h0;
  assign mem_MPORT_51_addr = 7'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 32'h0;
  assign mem_MPORT_52_addr = 7'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 32'h0;
  assign mem_MPORT_53_addr = 7'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 32'h0;
  assign mem_MPORT_54_addr = 7'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 32'h0;
  assign mem_MPORT_55_addr = 7'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 32'h0;
  assign mem_MPORT_56_addr = 7'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 32'h0;
  assign mem_MPORT_57_addr = 7'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 32'h0;
  assign mem_MPORT_58_addr = 7'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 32'h0;
  assign mem_MPORT_59_addr = 7'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 32'h0;
  assign mem_MPORT_60_addr = 7'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 32'h0;
  assign mem_MPORT_61_addr = 7'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 32'h0;
  assign mem_MPORT_62_addr = 7'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 32'h0;
  assign mem_MPORT_63_addr = 7'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 32'h0;
  assign mem_MPORT_64_addr = 7'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 32'h0;
  assign mem_MPORT_65_addr = 7'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 32'h0;
  assign mem_MPORT_66_addr = 7'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 32'h0;
  assign mem_MPORT_67_addr = 7'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 32'h0;
  assign mem_MPORT_68_addr = 7'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 32'h0;
  assign mem_MPORT_69_addr = 7'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 32'h0;
  assign mem_MPORT_70_addr = 7'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 32'h0;
  assign mem_MPORT_71_addr = 7'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 32'h0;
  assign mem_MPORT_72_addr = 7'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 32'h0;
  assign mem_MPORT_73_addr = 7'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 32'h0;
  assign mem_MPORT_74_addr = 7'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 32'h0;
  assign mem_MPORT_75_addr = 7'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 32'h0;
  assign mem_MPORT_76_addr = 7'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 32'h0;
  assign mem_MPORT_77_addr = 7'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 32'h0;
  assign mem_MPORT_78_addr = 7'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 32'h0;
  assign mem_MPORT_79_addr = 7'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 32'h0;
  assign mem_MPORT_80_addr = 7'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 32'h0;
  assign mem_MPORT_81_addr = 7'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 32'h0;
  assign mem_MPORT_82_addr = 7'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 32'h0;
  assign mem_MPORT_83_addr = 7'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 32'h0;
  assign mem_MPORT_84_addr = 7'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 32'h0;
  assign mem_MPORT_85_addr = 7'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 32'h0;
  assign mem_MPORT_86_addr = 7'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 32'h0;
  assign mem_MPORT_87_addr = 7'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 32'h0;
  assign mem_MPORT_88_addr = 7'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 32'h0;
  assign mem_MPORT_89_addr = 7'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 32'h0;
  assign mem_MPORT_90_addr = 7'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 32'h0;
  assign mem_MPORT_91_addr = 7'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 32'h0;
  assign mem_MPORT_92_addr = 7'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 32'h0;
  assign mem_MPORT_93_addr = 7'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 32'h0;
  assign mem_MPORT_94_addr = 7'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 32'h0;
  assign mem_MPORT_95_addr = 7'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 32'h0;
  assign mem_MPORT_96_addr = 7'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 32'h0;
  assign mem_MPORT_97_addr = 7'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 32'h0;
  assign mem_MPORT_98_addr = 7'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 32'h0;
  assign mem_MPORT_99_addr = 7'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 32'h0;
  assign mem_MPORT_100_addr = 7'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 32'h0;
  assign mem_MPORT_101_addr = 7'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 32'h0;
  assign mem_MPORT_102_addr = 7'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 32'h0;
  assign mem_MPORT_103_addr = 7'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 32'h0;
  assign mem_MPORT_104_addr = 7'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 32'h0;
  assign mem_MPORT_105_addr = 7'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 32'h0;
  assign mem_MPORT_106_addr = 7'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 32'h0;
  assign mem_MPORT_107_addr = 7'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 32'h0;
  assign mem_MPORT_108_addr = 7'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 32'h0;
  assign mem_MPORT_109_addr = 7'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 32'h0;
  assign mem_MPORT_110_addr = 7'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 32'h0;
  assign mem_MPORT_111_addr = 7'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 32'h0;
  assign mem_MPORT_112_addr = 7'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 32'h0;
  assign mem_MPORT_113_addr = 7'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 32'h0;
  assign mem_MPORT_114_addr = 7'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 32'h0;
  assign mem_MPORT_115_addr = 7'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 32'h0;
  assign mem_MPORT_116_addr = 7'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 32'h0;
  assign mem_MPORT_117_addr = 7'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 32'h0;
  assign mem_MPORT_118_addr = 7'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 32'h0;
  assign mem_MPORT_119_addr = 7'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 32'h0;
  assign mem_MPORT_120_addr = 7'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 32'h0;
  assign mem_MPORT_121_addr = 7'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 32'h0;
  assign mem_MPORT_122_addr = 7'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 32'h0;
  assign mem_MPORT_123_addr = 7'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 32'h0;
  assign mem_MPORT_124_addr = 7'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 32'h0;
  assign mem_MPORT_125_addr = 7'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 32'h0;
  assign mem_MPORT_126_addr = 7'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 32'h0;
  assign mem_MPORT_127_addr = 7'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = io_w_data;
  assign mem_MPORT_128_addr = io_w_addr;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P(
  input         clock,
  input         reset,
  input  [6:0]  io_r_addr,
  output [31:0] io_r_data_0,
  output [31:0] io_r_data_1,
  output [31:0] io_r_data_2,
  output [31:0] io_r_data_3,
  output [31:0] io_r_data_4,
  output [31:0] io_r_data_5,
  output [31:0] io_r_data_6,
  output [31:0] io_r_data_7,
  input         io_w_en,
  input  [6:0]  io_w_addr,
  input  [31:0] io_w_data_0,
  input  [31:0] io_w_data_1,
  input  [31:0] io_w_data_2,
  input  [31:0] io_w_data_3,
  input  [31:0] io_w_data_4,
  input  [31:0] io_w_data_5,
  input  [31:0] io_w_data_6,
  input  [31:0] io_w_data_7,
  input  [7:0]  io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_clock; // @[SRAM_1.scala 201:38]
  wire  brams_4_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_4_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_4_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_clock; // @[SRAM_1.scala 201:38]
  wire  brams_5_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_5_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_5_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_clock; // @[SRAM_1.scala 201:38]
  wire  brams_6_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_6_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_6_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_clock; // @[SRAM_1.scala 201:38]
  wire  brams_7_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_7_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_7_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  BankRAM_2P brams_4 ( // @[SRAM_1.scala 201:38]
    .clock(brams_4_clock),
    .reset(brams_4_reset),
    .io_r_addr(brams_4_io_r_addr),
    .io_r_data(brams_4_io_r_data),
    .io_w_en(brams_4_io_w_en),
    .io_w_addr(brams_4_io_w_addr),
    .io_w_data(brams_4_io_w_data)
  );
  BankRAM_2P brams_5 ( // @[SRAM_1.scala 201:38]
    .clock(brams_5_clock),
    .reset(brams_5_reset),
    .io_r_addr(brams_5_io_r_addr),
    .io_r_data(brams_5_io_r_data),
    .io_w_en(brams_5_io_w_en),
    .io_w_addr(brams_5_io_w_addr),
    .io_w_data(brams_5_io_w_data)
  );
  BankRAM_2P brams_6 ( // @[SRAM_1.scala 201:38]
    .clock(brams_6_clock),
    .reset(brams_6_reset),
    .io_r_addr(brams_6_io_r_addr),
    .io_r_data(brams_6_io_r_data),
    .io_w_en(brams_6_io_w_en),
    .io_w_addr(brams_6_io_w_addr),
    .io_w_data(brams_6_io_w_data)
  );
  BankRAM_2P brams_7 ( // @[SRAM_1.scala 201:38]
    .clock(brams_7_clock),
    .reset(brams_7_reset),
    .io_r_addr(brams_7_io_r_addr),
    .io_r_data(brams_7_io_r_data),
    .io_w_en(brams_7_io_w_en),
    .io_w_addr(brams_7_io_w_addr),
    .io_w_data(brams_7_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_4 = brams_4_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_5 = brams_5_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_6 = brams_6_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_7 = brams_7_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
  assign brams_4_clock = clock;
  assign brams_4_reset = reset;
  assign brams_4_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_4_io_w_en = io_w_en & io_w_maskOH[4]; // @[SRAM_1.scala 208:37]
  assign brams_4_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_4_io_w_data = io_w_data_4; // @[SRAM_1.scala 210:28]
  assign brams_5_clock = clock;
  assign brams_5_reset = reset;
  assign brams_5_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_5_io_w_en = io_w_en & io_w_maskOH[5]; // @[SRAM_1.scala 208:37]
  assign brams_5_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_5_io_w_data = io_w_data_5; // @[SRAM_1.scala 210:28]
  assign brams_6_clock = clock;
  assign brams_6_reset = reset;
  assign brams_6_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_6_io_w_en = io_w_en & io_w_maskOH[6]; // @[SRAM_1.scala 208:37]
  assign brams_6_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_6_io_w_data = io_w_data_6; // @[SRAM_1.scala 210:28]
  assign brams_7_clock = clock;
  assign brams_7_reset = reset;
  assign brams_7_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_7_io_w_en = io_w_en & io_w_maskOH[7]; // @[SRAM_1.scala 208:37]
  assign brams_7_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_7_io_w_data = io_w_data_7; // @[SRAM_1.scala 210:28]
endmodule
module DataBankArray(
  input         clock,
  input         reset,
  output        io_read_req_ready,
  input         io_read_req_valid,
  input  [6:0]  io_read_req_bits_set,
  output [31:0] io_read_resp_0_0,
  output [31:0] io_read_resp_0_1,
  output [31:0] io_read_resp_0_2,
  output [31:0] io_read_resp_0_3,
  output [31:0] io_read_resp_0_4,
  output [31:0] io_read_resp_0_5,
  output [31:0] io_read_resp_0_6,
  output [31:0] io_read_resp_0_7,
  output [31:0] io_read_resp_1_0,
  output [31:0] io_read_resp_1_1,
  output [31:0] io_read_resp_1_2,
  output [31:0] io_read_resp_1_3,
  output [31:0] io_read_resp_1_4,
  output [31:0] io_read_resp_1_5,
  output [31:0] io_read_resp_1_6,
  output [31:0] io_read_resp_1_7,
  output [31:0] io_read_resp_2_0,
  output [31:0] io_read_resp_2_1,
  output [31:0] io_read_resp_2_2,
  output [31:0] io_read_resp_2_3,
  output [31:0] io_read_resp_2_4,
  output [31:0] io_read_resp_2_5,
  output [31:0] io_read_resp_2_6,
  output [31:0] io_read_resp_2_7,
  output [31:0] io_read_resp_3_0,
  output [31:0] io_read_resp_3_1,
  output [31:0] io_read_resp_3_2,
  output [31:0] io_read_resp_3_3,
  output [31:0] io_read_resp_3_4,
  output [31:0] io_read_resp_3_5,
  output [31:0] io_read_resp_3_6,
  output [31:0] io_read_resp_3_7,
  output [31:0] io_read_resp_4_0,
  output [31:0] io_read_resp_4_1,
  output [31:0] io_read_resp_4_2,
  output [31:0] io_read_resp_4_3,
  output [31:0] io_read_resp_4_4,
  output [31:0] io_read_resp_4_5,
  output [31:0] io_read_resp_4_6,
  output [31:0] io_read_resp_4_7,
  output [31:0] io_read_resp_5_0,
  output [31:0] io_read_resp_5_1,
  output [31:0] io_read_resp_5_2,
  output [31:0] io_read_resp_5_3,
  output [31:0] io_read_resp_5_4,
  output [31:0] io_read_resp_5_5,
  output [31:0] io_read_resp_5_6,
  output [31:0] io_read_resp_5_7,
  output [31:0] io_read_resp_6_0,
  output [31:0] io_read_resp_6_1,
  output [31:0] io_read_resp_6_2,
  output [31:0] io_read_resp_6_3,
  output [31:0] io_read_resp_6_4,
  output [31:0] io_read_resp_6_5,
  output [31:0] io_read_resp_6_6,
  output [31:0] io_read_resp_6_7,
  output [31:0] io_read_resp_7_0,
  output [31:0] io_read_resp_7_1,
  output [31:0] io_read_resp_7_2,
  output [31:0] io_read_resp_7_3,
  output [31:0] io_read_resp_7_4,
  output [31:0] io_read_resp_7_5,
  output [31:0] io_read_resp_7_6,
  output [31:0] io_read_resp_7_7,
  output        io_write_req_ready,
  input         io_write_req_valid,
  input  [6:0]  io_write_req_bits_set,
  input  [31:0] io_write_req_bits_data_0,
  input  [31:0] io_write_req_bits_data_1,
  input  [31:0] io_write_req_bits_data_2,
  input  [31:0] io_write_req_bits_data_3,
  input  [31:0] io_write_req_bits_data_4,
  input  [31:0] io_write_req_bits_data_5,
  input  [31:0] io_write_req_bits_data_6,
  input  [31:0] io_write_req_bits_data_7,
  input  [7:0]  io_write_req_bits_blockMask,
  input  [7:0]  io_write_req_bits_way
);
  wire  dataBanks_0_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_0_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_0_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_0_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_0_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_0_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_1_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_1_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_1_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_2_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_2_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_2_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_3_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_3_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_3_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_4_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_4_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_4_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_4_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_4_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_4_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_5_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_5_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_5_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_5_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_5_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_5_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_6_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_6_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_6_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_6_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_6_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_6_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_7_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_7_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_7_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  dataBanks_7_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] dataBanks_7_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_7_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  ren = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  wire  _wen_T_1 = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  SRAMArray_2P dataBanks_0 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_0_clock),
    .reset(dataBanks_0_reset),
    .io_r_addr(dataBanks_0_io_r_addr),
    .io_r_data_0(dataBanks_0_io_r_data_0),
    .io_r_data_1(dataBanks_0_io_r_data_1),
    .io_r_data_2(dataBanks_0_io_r_data_2),
    .io_r_data_3(dataBanks_0_io_r_data_3),
    .io_r_data_4(dataBanks_0_io_r_data_4),
    .io_r_data_5(dataBanks_0_io_r_data_5),
    .io_r_data_6(dataBanks_0_io_r_data_6),
    .io_r_data_7(dataBanks_0_io_r_data_7),
    .io_w_en(dataBanks_0_io_w_en),
    .io_w_addr(dataBanks_0_io_w_addr),
    .io_w_data_0(dataBanks_0_io_w_data_0),
    .io_w_data_1(dataBanks_0_io_w_data_1),
    .io_w_data_2(dataBanks_0_io_w_data_2),
    .io_w_data_3(dataBanks_0_io_w_data_3),
    .io_w_data_4(dataBanks_0_io_w_data_4),
    .io_w_data_5(dataBanks_0_io_w_data_5),
    .io_w_data_6(dataBanks_0_io_w_data_6),
    .io_w_data_7(dataBanks_0_io_w_data_7),
    .io_w_maskOH(dataBanks_0_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_1 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_1_clock),
    .reset(dataBanks_1_reset),
    .io_r_addr(dataBanks_1_io_r_addr),
    .io_r_data_0(dataBanks_1_io_r_data_0),
    .io_r_data_1(dataBanks_1_io_r_data_1),
    .io_r_data_2(dataBanks_1_io_r_data_2),
    .io_r_data_3(dataBanks_1_io_r_data_3),
    .io_r_data_4(dataBanks_1_io_r_data_4),
    .io_r_data_5(dataBanks_1_io_r_data_5),
    .io_r_data_6(dataBanks_1_io_r_data_6),
    .io_r_data_7(dataBanks_1_io_r_data_7),
    .io_w_en(dataBanks_1_io_w_en),
    .io_w_addr(dataBanks_1_io_w_addr),
    .io_w_data_0(dataBanks_1_io_w_data_0),
    .io_w_data_1(dataBanks_1_io_w_data_1),
    .io_w_data_2(dataBanks_1_io_w_data_2),
    .io_w_data_3(dataBanks_1_io_w_data_3),
    .io_w_data_4(dataBanks_1_io_w_data_4),
    .io_w_data_5(dataBanks_1_io_w_data_5),
    .io_w_data_6(dataBanks_1_io_w_data_6),
    .io_w_data_7(dataBanks_1_io_w_data_7),
    .io_w_maskOH(dataBanks_1_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_2 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_2_clock),
    .reset(dataBanks_2_reset),
    .io_r_addr(dataBanks_2_io_r_addr),
    .io_r_data_0(dataBanks_2_io_r_data_0),
    .io_r_data_1(dataBanks_2_io_r_data_1),
    .io_r_data_2(dataBanks_2_io_r_data_2),
    .io_r_data_3(dataBanks_2_io_r_data_3),
    .io_r_data_4(dataBanks_2_io_r_data_4),
    .io_r_data_5(dataBanks_2_io_r_data_5),
    .io_r_data_6(dataBanks_2_io_r_data_6),
    .io_r_data_7(dataBanks_2_io_r_data_7),
    .io_w_en(dataBanks_2_io_w_en),
    .io_w_addr(dataBanks_2_io_w_addr),
    .io_w_data_0(dataBanks_2_io_w_data_0),
    .io_w_data_1(dataBanks_2_io_w_data_1),
    .io_w_data_2(dataBanks_2_io_w_data_2),
    .io_w_data_3(dataBanks_2_io_w_data_3),
    .io_w_data_4(dataBanks_2_io_w_data_4),
    .io_w_data_5(dataBanks_2_io_w_data_5),
    .io_w_data_6(dataBanks_2_io_w_data_6),
    .io_w_data_7(dataBanks_2_io_w_data_7),
    .io_w_maskOH(dataBanks_2_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_3 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_3_clock),
    .reset(dataBanks_3_reset),
    .io_r_addr(dataBanks_3_io_r_addr),
    .io_r_data_0(dataBanks_3_io_r_data_0),
    .io_r_data_1(dataBanks_3_io_r_data_1),
    .io_r_data_2(dataBanks_3_io_r_data_2),
    .io_r_data_3(dataBanks_3_io_r_data_3),
    .io_r_data_4(dataBanks_3_io_r_data_4),
    .io_r_data_5(dataBanks_3_io_r_data_5),
    .io_r_data_6(dataBanks_3_io_r_data_6),
    .io_r_data_7(dataBanks_3_io_r_data_7),
    .io_w_en(dataBanks_3_io_w_en),
    .io_w_addr(dataBanks_3_io_w_addr),
    .io_w_data_0(dataBanks_3_io_w_data_0),
    .io_w_data_1(dataBanks_3_io_w_data_1),
    .io_w_data_2(dataBanks_3_io_w_data_2),
    .io_w_data_3(dataBanks_3_io_w_data_3),
    .io_w_data_4(dataBanks_3_io_w_data_4),
    .io_w_data_5(dataBanks_3_io_w_data_5),
    .io_w_data_6(dataBanks_3_io_w_data_6),
    .io_w_data_7(dataBanks_3_io_w_data_7),
    .io_w_maskOH(dataBanks_3_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_4 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_4_clock),
    .reset(dataBanks_4_reset),
    .io_r_addr(dataBanks_4_io_r_addr),
    .io_r_data_0(dataBanks_4_io_r_data_0),
    .io_r_data_1(dataBanks_4_io_r_data_1),
    .io_r_data_2(dataBanks_4_io_r_data_2),
    .io_r_data_3(dataBanks_4_io_r_data_3),
    .io_r_data_4(dataBanks_4_io_r_data_4),
    .io_r_data_5(dataBanks_4_io_r_data_5),
    .io_r_data_6(dataBanks_4_io_r_data_6),
    .io_r_data_7(dataBanks_4_io_r_data_7),
    .io_w_en(dataBanks_4_io_w_en),
    .io_w_addr(dataBanks_4_io_w_addr),
    .io_w_data_0(dataBanks_4_io_w_data_0),
    .io_w_data_1(dataBanks_4_io_w_data_1),
    .io_w_data_2(dataBanks_4_io_w_data_2),
    .io_w_data_3(dataBanks_4_io_w_data_3),
    .io_w_data_4(dataBanks_4_io_w_data_4),
    .io_w_data_5(dataBanks_4_io_w_data_5),
    .io_w_data_6(dataBanks_4_io_w_data_6),
    .io_w_data_7(dataBanks_4_io_w_data_7),
    .io_w_maskOH(dataBanks_4_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_5 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_5_clock),
    .reset(dataBanks_5_reset),
    .io_r_addr(dataBanks_5_io_r_addr),
    .io_r_data_0(dataBanks_5_io_r_data_0),
    .io_r_data_1(dataBanks_5_io_r_data_1),
    .io_r_data_2(dataBanks_5_io_r_data_2),
    .io_r_data_3(dataBanks_5_io_r_data_3),
    .io_r_data_4(dataBanks_5_io_r_data_4),
    .io_r_data_5(dataBanks_5_io_r_data_5),
    .io_r_data_6(dataBanks_5_io_r_data_6),
    .io_r_data_7(dataBanks_5_io_r_data_7),
    .io_w_en(dataBanks_5_io_w_en),
    .io_w_addr(dataBanks_5_io_w_addr),
    .io_w_data_0(dataBanks_5_io_w_data_0),
    .io_w_data_1(dataBanks_5_io_w_data_1),
    .io_w_data_2(dataBanks_5_io_w_data_2),
    .io_w_data_3(dataBanks_5_io_w_data_3),
    .io_w_data_4(dataBanks_5_io_w_data_4),
    .io_w_data_5(dataBanks_5_io_w_data_5),
    .io_w_data_6(dataBanks_5_io_w_data_6),
    .io_w_data_7(dataBanks_5_io_w_data_7),
    .io_w_maskOH(dataBanks_5_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_6 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_6_clock),
    .reset(dataBanks_6_reset),
    .io_r_addr(dataBanks_6_io_r_addr),
    .io_r_data_0(dataBanks_6_io_r_data_0),
    .io_r_data_1(dataBanks_6_io_r_data_1),
    .io_r_data_2(dataBanks_6_io_r_data_2),
    .io_r_data_3(dataBanks_6_io_r_data_3),
    .io_r_data_4(dataBanks_6_io_r_data_4),
    .io_r_data_5(dataBanks_6_io_r_data_5),
    .io_r_data_6(dataBanks_6_io_r_data_6),
    .io_r_data_7(dataBanks_6_io_r_data_7),
    .io_w_en(dataBanks_6_io_w_en),
    .io_w_addr(dataBanks_6_io_w_addr),
    .io_w_data_0(dataBanks_6_io_w_data_0),
    .io_w_data_1(dataBanks_6_io_w_data_1),
    .io_w_data_2(dataBanks_6_io_w_data_2),
    .io_w_data_3(dataBanks_6_io_w_data_3),
    .io_w_data_4(dataBanks_6_io_w_data_4),
    .io_w_data_5(dataBanks_6_io_w_data_5),
    .io_w_data_6(dataBanks_6_io_w_data_6),
    .io_w_data_7(dataBanks_6_io_w_data_7),
    .io_w_maskOH(dataBanks_6_io_w_maskOH)
  );
  SRAMArray_2P dataBanks_7 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_7_clock),
    .reset(dataBanks_7_reset),
    .io_r_addr(dataBanks_7_io_r_addr),
    .io_r_data_0(dataBanks_7_io_r_data_0),
    .io_r_data_1(dataBanks_7_io_r_data_1),
    .io_r_data_2(dataBanks_7_io_r_data_2),
    .io_r_data_3(dataBanks_7_io_r_data_3),
    .io_r_data_4(dataBanks_7_io_r_data_4),
    .io_r_data_5(dataBanks_7_io_r_data_5),
    .io_r_data_6(dataBanks_7_io_r_data_6),
    .io_r_data_7(dataBanks_7_io_r_data_7),
    .io_w_en(dataBanks_7_io_w_en),
    .io_w_addr(dataBanks_7_io_w_addr),
    .io_w_data_0(dataBanks_7_io_w_data_0),
    .io_w_data_1(dataBanks_7_io_w_data_1),
    .io_w_data_2(dataBanks_7_io_w_data_2),
    .io_w_data_3(dataBanks_7_io_w_data_3),
    .io_w_data_4(dataBanks_7_io_w_data_4),
    .io_w_data_5(dataBanks_7_io_w_data_5),
    .io_w_data_6(dataBanks_7_io_w_data_6),
    .io_w_data_7(dataBanks_7_io_w_data_7),
    .io_w_maskOH(dataBanks_7_io_w_maskOH)
  );
  assign io_read_req_ready = 1'h1; // @[DataBank.scala 46:23]
  assign io_read_resp_0_0 = ren ? dataBanks_0_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_1 = ren ? dataBanks_0_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_2 = ren ? dataBanks_0_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_3 = ren ? dataBanks_0_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_4 = ren ? dataBanks_0_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_5 = ren ? dataBanks_0_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_6 = ren ? dataBanks_0_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_7 = ren ? dataBanks_0_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_0 = ren ? dataBanks_1_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_1 = ren ? dataBanks_1_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_2 = ren ? dataBanks_1_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_3 = ren ? dataBanks_1_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_4 = ren ? dataBanks_1_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_5 = ren ? dataBanks_1_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_6 = ren ? dataBanks_1_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_7 = ren ? dataBanks_1_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_0 = ren ? dataBanks_2_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_1 = ren ? dataBanks_2_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_2 = ren ? dataBanks_2_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_3 = ren ? dataBanks_2_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_4 = ren ? dataBanks_2_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_5 = ren ? dataBanks_2_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_6 = ren ? dataBanks_2_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_7 = ren ? dataBanks_2_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_0 = ren ? dataBanks_3_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_1 = ren ? dataBanks_3_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_2 = ren ? dataBanks_3_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_3 = ren ? dataBanks_3_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_4 = ren ? dataBanks_3_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_5 = ren ? dataBanks_3_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_6 = ren ? dataBanks_3_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_7 = ren ? dataBanks_3_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_0 = ren ? dataBanks_4_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_1 = ren ? dataBanks_4_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_2 = ren ? dataBanks_4_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_3 = ren ? dataBanks_4_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_4 = ren ? dataBanks_4_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_5 = ren ? dataBanks_4_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_6 = ren ? dataBanks_4_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_7 = ren ? dataBanks_4_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_0 = ren ? dataBanks_5_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_1 = ren ? dataBanks_5_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_2 = ren ? dataBanks_5_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_3 = ren ? dataBanks_5_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_4 = ren ? dataBanks_5_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_5 = ren ? dataBanks_5_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_6 = ren ? dataBanks_5_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_7 = ren ? dataBanks_5_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_0 = ren ? dataBanks_6_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_1 = ren ? dataBanks_6_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_2 = ren ? dataBanks_6_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_3 = ren ? dataBanks_6_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_4 = ren ? dataBanks_6_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_5 = ren ? dataBanks_6_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_6 = ren ? dataBanks_6_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_7 = ren ? dataBanks_6_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_0 = ren ? dataBanks_7_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_1 = ren ? dataBanks_7_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_2 = ren ? dataBanks_7_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_3 = ren ? dataBanks_7_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_4 = ren ? dataBanks_7_io_r_data_4 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_5 = ren ? dataBanks_7_io_r_data_5 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_6 = ren ? dataBanks_7_io_r_data_6 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_7 = ren ? dataBanks_7_io_r_data_7 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_write_req_ready = 1'h1; // @[DataBank.scala 55:28]
  assign dataBanks_0_clock = clock;
  assign dataBanks_0_reset = reset;
  assign dataBanks_0_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_0_io_w_en = io_write_req_bits_way[0] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_0_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_0_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_1_clock = clock;
  assign dataBanks_1_reset = reset;
  assign dataBanks_1_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_1_io_w_en = io_write_req_bits_way[1] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_1_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_1_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_2_clock = clock;
  assign dataBanks_2_reset = reset;
  assign dataBanks_2_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_2_io_w_en = io_write_req_bits_way[2] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_2_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_2_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_3_clock = clock;
  assign dataBanks_3_reset = reset;
  assign dataBanks_3_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_3_io_w_en = io_write_req_bits_way[3] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_3_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_3_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_4_clock = clock;
  assign dataBanks_4_reset = reset;
  assign dataBanks_4_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_4_io_w_en = io_write_req_bits_way[4] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_4_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_4_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_5_clock = clock;
  assign dataBanks_5_reset = reset;
  assign dataBanks_5_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_5_io_w_en = io_write_req_bits_way[5] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_5_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_5_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_6_clock = clock;
  assign dataBanks_6_reset = reset;
  assign dataBanks_6_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_6_io_w_en = io_write_req_bits_way[6] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_6_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_6_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_7_clock = clock;
  assign dataBanks_7_reset = reset;
  assign dataBanks_7_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_7_io_w_en = io_write_req_bits_way[7] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_7_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_7_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_4 = io_write_req_bits_data_4; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_5 = io_write_req_bits_data_5; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_6 = io_write_req_bits_data_6; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_7 = io_write_req_bits_data_7; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
endmodule
module BankRAM_2P_64(
  input         clock,
  input         reset,
  input  [6:0]  io_r_addr,
  output [19:0] io_r_data,
  input         io_w_en,
  input  [6:0]  io_w_addr,
  input  [19:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] mem [0:127]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [6:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 20'h0;
  assign mem_MPORT_addr = 7'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 20'h0;
  assign mem_MPORT_1_addr = 7'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 20'h0;
  assign mem_MPORT_2_addr = 7'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 20'h0;
  assign mem_MPORT_3_addr = 7'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 20'h0;
  assign mem_MPORT_4_addr = 7'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 20'h0;
  assign mem_MPORT_5_addr = 7'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 20'h0;
  assign mem_MPORT_6_addr = 7'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 20'h0;
  assign mem_MPORT_7_addr = 7'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 20'h0;
  assign mem_MPORT_8_addr = 7'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 20'h0;
  assign mem_MPORT_9_addr = 7'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 20'h0;
  assign mem_MPORT_10_addr = 7'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 20'h0;
  assign mem_MPORT_11_addr = 7'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 20'h0;
  assign mem_MPORT_12_addr = 7'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 20'h0;
  assign mem_MPORT_13_addr = 7'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 20'h0;
  assign mem_MPORT_14_addr = 7'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 20'h0;
  assign mem_MPORT_15_addr = 7'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 20'h0;
  assign mem_MPORT_16_addr = 7'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 20'h0;
  assign mem_MPORT_17_addr = 7'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 20'h0;
  assign mem_MPORT_18_addr = 7'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 20'h0;
  assign mem_MPORT_19_addr = 7'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 20'h0;
  assign mem_MPORT_20_addr = 7'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 20'h0;
  assign mem_MPORT_21_addr = 7'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 20'h0;
  assign mem_MPORT_22_addr = 7'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 20'h0;
  assign mem_MPORT_23_addr = 7'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 20'h0;
  assign mem_MPORT_24_addr = 7'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 20'h0;
  assign mem_MPORT_25_addr = 7'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 20'h0;
  assign mem_MPORT_26_addr = 7'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 20'h0;
  assign mem_MPORT_27_addr = 7'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 20'h0;
  assign mem_MPORT_28_addr = 7'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 20'h0;
  assign mem_MPORT_29_addr = 7'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 20'h0;
  assign mem_MPORT_30_addr = 7'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 20'h0;
  assign mem_MPORT_31_addr = 7'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 20'h0;
  assign mem_MPORT_32_addr = 7'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 20'h0;
  assign mem_MPORT_33_addr = 7'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 20'h0;
  assign mem_MPORT_34_addr = 7'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 20'h0;
  assign mem_MPORT_35_addr = 7'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 20'h0;
  assign mem_MPORT_36_addr = 7'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 20'h0;
  assign mem_MPORT_37_addr = 7'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 20'h0;
  assign mem_MPORT_38_addr = 7'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 20'h0;
  assign mem_MPORT_39_addr = 7'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 20'h0;
  assign mem_MPORT_40_addr = 7'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 20'h0;
  assign mem_MPORT_41_addr = 7'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 20'h0;
  assign mem_MPORT_42_addr = 7'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 20'h0;
  assign mem_MPORT_43_addr = 7'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 20'h0;
  assign mem_MPORT_44_addr = 7'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 20'h0;
  assign mem_MPORT_45_addr = 7'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 20'h0;
  assign mem_MPORT_46_addr = 7'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 20'h0;
  assign mem_MPORT_47_addr = 7'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 20'h0;
  assign mem_MPORT_48_addr = 7'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 20'h0;
  assign mem_MPORT_49_addr = 7'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 20'h0;
  assign mem_MPORT_50_addr = 7'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 20'h0;
  assign mem_MPORT_51_addr = 7'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 20'h0;
  assign mem_MPORT_52_addr = 7'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 20'h0;
  assign mem_MPORT_53_addr = 7'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 20'h0;
  assign mem_MPORT_54_addr = 7'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 20'h0;
  assign mem_MPORT_55_addr = 7'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 20'h0;
  assign mem_MPORT_56_addr = 7'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 20'h0;
  assign mem_MPORT_57_addr = 7'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 20'h0;
  assign mem_MPORT_58_addr = 7'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 20'h0;
  assign mem_MPORT_59_addr = 7'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 20'h0;
  assign mem_MPORT_60_addr = 7'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 20'h0;
  assign mem_MPORT_61_addr = 7'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 20'h0;
  assign mem_MPORT_62_addr = 7'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 20'h0;
  assign mem_MPORT_63_addr = 7'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 20'h0;
  assign mem_MPORT_64_addr = 7'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 20'h0;
  assign mem_MPORT_65_addr = 7'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 20'h0;
  assign mem_MPORT_66_addr = 7'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 20'h0;
  assign mem_MPORT_67_addr = 7'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 20'h0;
  assign mem_MPORT_68_addr = 7'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 20'h0;
  assign mem_MPORT_69_addr = 7'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 20'h0;
  assign mem_MPORT_70_addr = 7'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 20'h0;
  assign mem_MPORT_71_addr = 7'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 20'h0;
  assign mem_MPORT_72_addr = 7'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 20'h0;
  assign mem_MPORT_73_addr = 7'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 20'h0;
  assign mem_MPORT_74_addr = 7'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 20'h0;
  assign mem_MPORT_75_addr = 7'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 20'h0;
  assign mem_MPORT_76_addr = 7'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 20'h0;
  assign mem_MPORT_77_addr = 7'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 20'h0;
  assign mem_MPORT_78_addr = 7'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 20'h0;
  assign mem_MPORT_79_addr = 7'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 20'h0;
  assign mem_MPORT_80_addr = 7'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 20'h0;
  assign mem_MPORT_81_addr = 7'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 20'h0;
  assign mem_MPORT_82_addr = 7'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 20'h0;
  assign mem_MPORT_83_addr = 7'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 20'h0;
  assign mem_MPORT_84_addr = 7'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 20'h0;
  assign mem_MPORT_85_addr = 7'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 20'h0;
  assign mem_MPORT_86_addr = 7'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 20'h0;
  assign mem_MPORT_87_addr = 7'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 20'h0;
  assign mem_MPORT_88_addr = 7'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 20'h0;
  assign mem_MPORT_89_addr = 7'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 20'h0;
  assign mem_MPORT_90_addr = 7'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 20'h0;
  assign mem_MPORT_91_addr = 7'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 20'h0;
  assign mem_MPORT_92_addr = 7'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 20'h0;
  assign mem_MPORT_93_addr = 7'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 20'h0;
  assign mem_MPORT_94_addr = 7'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 20'h0;
  assign mem_MPORT_95_addr = 7'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 20'h0;
  assign mem_MPORT_96_addr = 7'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 20'h0;
  assign mem_MPORT_97_addr = 7'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 20'h0;
  assign mem_MPORT_98_addr = 7'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 20'h0;
  assign mem_MPORT_99_addr = 7'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 20'h0;
  assign mem_MPORT_100_addr = 7'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 20'h0;
  assign mem_MPORT_101_addr = 7'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 20'h0;
  assign mem_MPORT_102_addr = 7'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 20'h0;
  assign mem_MPORT_103_addr = 7'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 20'h0;
  assign mem_MPORT_104_addr = 7'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 20'h0;
  assign mem_MPORT_105_addr = 7'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 20'h0;
  assign mem_MPORT_106_addr = 7'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 20'h0;
  assign mem_MPORT_107_addr = 7'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 20'h0;
  assign mem_MPORT_108_addr = 7'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 20'h0;
  assign mem_MPORT_109_addr = 7'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 20'h0;
  assign mem_MPORT_110_addr = 7'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 20'h0;
  assign mem_MPORT_111_addr = 7'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 20'h0;
  assign mem_MPORT_112_addr = 7'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 20'h0;
  assign mem_MPORT_113_addr = 7'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 20'h0;
  assign mem_MPORT_114_addr = 7'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 20'h0;
  assign mem_MPORT_115_addr = 7'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 20'h0;
  assign mem_MPORT_116_addr = 7'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 20'h0;
  assign mem_MPORT_117_addr = 7'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 20'h0;
  assign mem_MPORT_118_addr = 7'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 20'h0;
  assign mem_MPORT_119_addr = 7'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 20'h0;
  assign mem_MPORT_120_addr = 7'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 20'h0;
  assign mem_MPORT_121_addr = 7'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 20'h0;
  assign mem_MPORT_122_addr = 7'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 20'h0;
  assign mem_MPORT_123_addr = 7'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 20'h0;
  assign mem_MPORT_124_addr = 7'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 20'h0;
  assign mem_MPORT_125_addr = 7'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 20'h0;
  assign mem_MPORT_126_addr = 7'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 20'h0;
  assign mem_MPORT_127_addr = 7'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = io_w_data;
  assign mem_MPORT_128_addr = io_w_addr;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_8(
  input         clock,
  input         reset,
  input  [6:0]  io_r_addr,
  output [19:0] io_r_data_0,
  output [19:0] io_r_data_1,
  output [19:0] io_r_data_2,
  output [19:0] io_r_data_3,
  output [19:0] io_r_data_4,
  output [19:0] io_r_data_5,
  output [19:0] io_r_data_6,
  output [19:0] io_r_data_7,
  input         io_w_en,
  input  [6:0]  io_w_addr,
  input  [19:0] io_w_data_0,
  input  [19:0] io_w_data_1,
  input  [19:0] io_w_data_2,
  input  [19:0] io_w_data_3,
  input  [19:0] io_w_data_4,
  input  [19:0] io_w_data_5,
  input  [19:0] io_w_data_6,
  input  [19:0] io_w_data_7,
  input  [7:0]  io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_clock; // @[SRAM_1.scala 201:38]
  wire  brams_4_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_4_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_4_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_clock; // @[SRAM_1.scala 201:38]
  wire  brams_5_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_5_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_5_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_clock; // @[SRAM_1.scala 201:38]
  wire  brams_6_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_6_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_6_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_clock; // @[SRAM_1.scala 201:38]
  wire  brams_7_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_7_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_7_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P_64 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P_64 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P_64 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P_64 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  BankRAM_2P_64 brams_4 ( // @[SRAM_1.scala 201:38]
    .clock(brams_4_clock),
    .reset(brams_4_reset),
    .io_r_addr(brams_4_io_r_addr),
    .io_r_data(brams_4_io_r_data),
    .io_w_en(brams_4_io_w_en),
    .io_w_addr(brams_4_io_w_addr),
    .io_w_data(brams_4_io_w_data)
  );
  BankRAM_2P_64 brams_5 ( // @[SRAM_1.scala 201:38]
    .clock(brams_5_clock),
    .reset(brams_5_reset),
    .io_r_addr(brams_5_io_r_addr),
    .io_r_data(brams_5_io_r_data),
    .io_w_en(brams_5_io_w_en),
    .io_w_addr(brams_5_io_w_addr),
    .io_w_data(brams_5_io_w_data)
  );
  BankRAM_2P_64 brams_6 ( // @[SRAM_1.scala 201:38]
    .clock(brams_6_clock),
    .reset(brams_6_reset),
    .io_r_addr(brams_6_io_r_addr),
    .io_r_data(brams_6_io_r_data),
    .io_w_en(brams_6_io_w_en),
    .io_w_addr(brams_6_io_w_addr),
    .io_w_data(brams_6_io_w_data)
  );
  BankRAM_2P_64 brams_7 ( // @[SRAM_1.scala 201:38]
    .clock(brams_7_clock),
    .reset(brams_7_reset),
    .io_r_addr(brams_7_io_r_addr),
    .io_r_data(brams_7_io_r_data),
    .io_w_en(brams_7_io_w_en),
    .io_w_addr(brams_7_io_w_addr),
    .io_w_data(brams_7_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_4 = brams_4_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_5 = brams_5_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_6 = brams_6_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_7 = brams_7_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
  assign brams_4_clock = clock;
  assign brams_4_reset = reset;
  assign brams_4_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_4_io_w_en = io_w_en & io_w_maskOH[4]; // @[SRAM_1.scala 208:37]
  assign brams_4_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_4_io_w_data = io_w_data_4; // @[SRAM_1.scala 210:28]
  assign brams_5_clock = clock;
  assign brams_5_reset = reset;
  assign brams_5_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_5_io_w_en = io_w_en & io_w_maskOH[5]; // @[SRAM_1.scala 208:37]
  assign brams_5_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_5_io_w_data = io_w_data_5; // @[SRAM_1.scala 210:28]
  assign brams_6_clock = clock;
  assign brams_6_reset = reset;
  assign brams_6_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_6_io_w_en = io_w_en & io_w_maskOH[6]; // @[SRAM_1.scala 208:37]
  assign brams_6_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_6_io_w_data = io_w_data_6; // @[SRAM_1.scala 210:28]
  assign brams_7_clock = clock;
  assign brams_7_reset = reset;
  assign brams_7_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_7_io_w_en = io_w_en & io_w_maskOH[7]; // @[SRAM_1.scala 208:37]
  assign brams_7_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_7_io_w_data = io_w_data_7; // @[SRAM_1.scala 210:28]
endmodule
module BankRAM_2P_72(
  input        clock,
  input        reset,
  input  [6:0] io_r_addr,
  output [1:0] io_r_data,
  input        io_w_en,
  input  [6:0] io_w_addr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] mem [0:127]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [6:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [6:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 2'h0;
  assign mem_MPORT_addr = 7'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 2'h0;
  assign mem_MPORT_1_addr = 7'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 2'h0;
  assign mem_MPORT_2_addr = 7'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 2'h0;
  assign mem_MPORT_3_addr = 7'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 2'h0;
  assign mem_MPORT_4_addr = 7'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 2'h0;
  assign mem_MPORT_5_addr = 7'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 2'h0;
  assign mem_MPORT_6_addr = 7'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 2'h0;
  assign mem_MPORT_7_addr = 7'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 2'h0;
  assign mem_MPORT_8_addr = 7'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 2'h0;
  assign mem_MPORT_9_addr = 7'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 2'h0;
  assign mem_MPORT_10_addr = 7'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 2'h0;
  assign mem_MPORT_11_addr = 7'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 2'h0;
  assign mem_MPORT_12_addr = 7'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 2'h0;
  assign mem_MPORT_13_addr = 7'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 2'h0;
  assign mem_MPORT_14_addr = 7'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 2'h0;
  assign mem_MPORT_15_addr = 7'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 2'h0;
  assign mem_MPORT_16_addr = 7'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 2'h0;
  assign mem_MPORT_17_addr = 7'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 2'h0;
  assign mem_MPORT_18_addr = 7'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 2'h0;
  assign mem_MPORT_19_addr = 7'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 2'h0;
  assign mem_MPORT_20_addr = 7'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 2'h0;
  assign mem_MPORT_21_addr = 7'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 2'h0;
  assign mem_MPORT_22_addr = 7'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 2'h0;
  assign mem_MPORT_23_addr = 7'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 2'h0;
  assign mem_MPORT_24_addr = 7'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 2'h0;
  assign mem_MPORT_25_addr = 7'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 2'h0;
  assign mem_MPORT_26_addr = 7'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 2'h0;
  assign mem_MPORT_27_addr = 7'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 2'h0;
  assign mem_MPORT_28_addr = 7'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 2'h0;
  assign mem_MPORT_29_addr = 7'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 2'h0;
  assign mem_MPORT_30_addr = 7'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 2'h0;
  assign mem_MPORT_31_addr = 7'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 2'h0;
  assign mem_MPORT_32_addr = 7'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 2'h0;
  assign mem_MPORT_33_addr = 7'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 2'h0;
  assign mem_MPORT_34_addr = 7'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 2'h0;
  assign mem_MPORT_35_addr = 7'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 2'h0;
  assign mem_MPORT_36_addr = 7'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 2'h0;
  assign mem_MPORT_37_addr = 7'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 2'h0;
  assign mem_MPORT_38_addr = 7'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 2'h0;
  assign mem_MPORT_39_addr = 7'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 2'h0;
  assign mem_MPORT_40_addr = 7'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 2'h0;
  assign mem_MPORT_41_addr = 7'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 2'h0;
  assign mem_MPORT_42_addr = 7'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 2'h0;
  assign mem_MPORT_43_addr = 7'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 2'h0;
  assign mem_MPORT_44_addr = 7'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 2'h0;
  assign mem_MPORT_45_addr = 7'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 2'h0;
  assign mem_MPORT_46_addr = 7'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 2'h0;
  assign mem_MPORT_47_addr = 7'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 2'h0;
  assign mem_MPORT_48_addr = 7'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 2'h0;
  assign mem_MPORT_49_addr = 7'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 2'h0;
  assign mem_MPORT_50_addr = 7'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 2'h0;
  assign mem_MPORT_51_addr = 7'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 2'h0;
  assign mem_MPORT_52_addr = 7'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 2'h0;
  assign mem_MPORT_53_addr = 7'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 2'h0;
  assign mem_MPORT_54_addr = 7'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 2'h0;
  assign mem_MPORT_55_addr = 7'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 2'h0;
  assign mem_MPORT_56_addr = 7'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 2'h0;
  assign mem_MPORT_57_addr = 7'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 2'h0;
  assign mem_MPORT_58_addr = 7'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 2'h0;
  assign mem_MPORT_59_addr = 7'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 2'h0;
  assign mem_MPORT_60_addr = 7'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 2'h0;
  assign mem_MPORT_61_addr = 7'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 2'h0;
  assign mem_MPORT_62_addr = 7'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 2'h0;
  assign mem_MPORT_63_addr = 7'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 2'h0;
  assign mem_MPORT_64_addr = 7'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 2'h0;
  assign mem_MPORT_65_addr = 7'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 2'h0;
  assign mem_MPORT_66_addr = 7'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 2'h0;
  assign mem_MPORT_67_addr = 7'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 2'h0;
  assign mem_MPORT_68_addr = 7'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 2'h0;
  assign mem_MPORT_69_addr = 7'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 2'h0;
  assign mem_MPORT_70_addr = 7'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 2'h0;
  assign mem_MPORT_71_addr = 7'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 2'h0;
  assign mem_MPORT_72_addr = 7'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 2'h0;
  assign mem_MPORT_73_addr = 7'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 2'h0;
  assign mem_MPORT_74_addr = 7'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 2'h0;
  assign mem_MPORT_75_addr = 7'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 2'h0;
  assign mem_MPORT_76_addr = 7'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 2'h0;
  assign mem_MPORT_77_addr = 7'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 2'h0;
  assign mem_MPORT_78_addr = 7'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 2'h0;
  assign mem_MPORT_79_addr = 7'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 2'h0;
  assign mem_MPORT_80_addr = 7'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 2'h0;
  assign mem_MPORT_81_addr = 7'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 2'h0;
  assign mem_MPORT_82_addr = 7'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 2'h0;
  assign mem_MPORT_83_addr = 7'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 2'h0;
  assign mem_MPORT_84_addr = 7'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 2'h0;
  assign mem_MPORT_85_addr = 7'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 2'h0;
  assign mem_MPORT_86_addr = 7'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 2'h0;
  assign mem_MPORT_87_addr = 7'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 2'h0;
  assign mem_MPORT_88_addr = 7'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 2'h0;
  assign mem_MPORT_89_addr = 7'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 2'h0;
  assign mem_MPORT_90_addr = 7'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 2'h0;
  assign mem_MPORT_91_addr = 7'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 2'h0;
  assign mem_MPORT_92_addr = 7'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 2'h0;
  assign mem_MPORT_93_addr = 7'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 2'h0;
  assign mem_MPORT_94_addr = 7'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 2'h0;
  assign mem_MPORT_95_addr = 7'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 2'h0;
  assign mem_MPORT_96_addr = 7'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 2'h0;
  assign mem_MPORT_97_addr = 7'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 2'h0;
  assign mem_MPORT_98_addr = 7'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 2'h0;
  assign mem_MPORT_99_addr = 7'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 2'h0;
  assign mem_MPORT_100_addr = 7'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 2'h0;
  assign mem_MPORT_101_addr = 7'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 2'h0;
  assign mem_MPORT_102_addr = 7'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 2'h0;
  assign mem_MPORT_103_addr = 7'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 2'h0;
  assign mem_MPORT_104_addr = 7'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 2'h0;
  assign mem_MPORT_105_addr = 7'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 2'h0;
  assign mem_MPORT_106_addr = 7'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 2'h0;
  assign mem_MPORT_107_addr = 7'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 2'h0;
  assign mem_MPORT_108_addr = 7'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 2'h0;
  assign mem_MPORT_109_addr = 7'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 2'h0;
  assign mem_MPORT_110_addr = 7'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 2'h0;
  assign mem_MPORT_111_addr = 7'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 2'h0;
  assign mem_MPORT_112_addr = 7'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 2'h0;
  assign mem_MPORT_113_addr = 7'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 2'h0;
  assign mem_MPORT_114_addr = 7'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 2'h0;
  assign mem_MPORT_115_addr = 7'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 2'h0;
  assign mem_MPORT_116_addr = 7'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 2'h0;
  assign mem_MPORT_117_addr = 7'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 2'h0;
  assign mem_MPORT_118_addr = 7'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 2'h0;
  assign mem_MPORT_119_addr = 7'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 2'h0;
  assign mem_MPORT_120_addr = 7'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 2'h0;
  assign mem_MPORT_121_addr = 7'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 2'h0;
  assign mem_MPORT_122_addr = 7'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 2'h0;
  assign mem_MPORT_123_addr = 7'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 2'h0;
  assign mem_MPORT_124_addr = 7'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 2'h0;
  assign mem_MPORT_125_addr = 7'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 2'h0;
  assign mem_MPORT_126_addr = 7'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 2'h0;
  assign mem_MPORT_127_addr = 7'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 2'h1;
  assign mem_MPORT_128_addr = io_w_addr;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? 2'h1 : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_9(
  input        clock,
  input        reset,
  input  [6:0] io_r_addr,
  output [1:0] io_r_data_0,
  output [1:0] io_r_data_1,
  output [1:0] io_r_data_2,
  output [1:0] io_r_data_3,
  output [1:0] io_r_data_4,
  output [1:0] io_r_data_5,
  output [1:0] io_r_data_6,
  output [1:0] io_r_data_7,
  input        io_w_en,
  input  [6:0] io_w_addr,
  input  [7:0] io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_4_clock; // @[SRAM_1.scala 201:38]
  wire  brams_4_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_4_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_4_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_5_clock; // @[SRAM_1.scala 201:38]
  wire  brams_5_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_5_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_5_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_6_clock; // @[SRAM_1.scala 201:38]
  wire  brams_6_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_6_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_6_io_w_addr; // @[SRAM_1.scala 201:38]
  wire  brams_7_clock; // @[SRAM_1.scala 201:38]
  wire  brams_7_reset; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_7_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_io_w_en; // @[SRAM_1.scala 201:38]
  wire [6:0] brams_7_io_w_addr; // @[SRAM_1.scala 201:38]
  BankRAM_2P_72 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr)
  );
  BankRAM_2P_72 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr)
  );
  BankRAM_2P_72 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr)
  );
  BankRAM_2P_72 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr)
  );
  BankRAM_2P_72 brams_4 ( // @[SRAM_1.scala 201:38]
    .clock(brams_4_clock),
    .reset(brams_4_reset),
    .io_r_addr(brams_4_io_r_addr),
    .io_r_data(brams_4_io_r_data),
    .io_w_en(brams_4_io_w_en),
    .io_w_addr(brams_4_io_w_addr)
  );
  BankRAM_2P_72 brams_5 ( // @[SRAM_1.scala 201:38]
    .clock(brams_5_clock),
    .reset(brams_5_reset),
    .io_r_addr(brams_5_io_r_addr),
    .io_r_data(brams_5_io_r_data),
    .io_w_en(brams_5_io_w_en),
    .io_w_addr(brams_5_io_w_addr)
  );
  BankRAM_2P_72 brams_6 ( // @[SRAM_1.scala 201:38]
    .clock(brams_6_clock),
    .reset(brams_6_reset),
    .io_r_addr(brams_6_io_r_addr),
    .io_r_data(brams_6_io_r_data),
    .io_w_en(brams_6_io_w_en),
    .io_w_addr(brams_6_io_w_addr)
  );
  BankRAM_2P_72 brams_7 ( // @[SRAM_1.scala 201:38]
    .clock(brams_7_clock),
    .reset(brams_7_reset),
    .io_r_addr(brams_7_io_r_addr),
    .io_r_data(brams_7_io_r_data),
    .io_w_en(brams_7_io_w_en),
    .io_w_addr(brams_7_io_w_addr)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_4 = brams_4_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_5 = brams_5_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_6 = brams_6_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_7 = brams_7_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_4_clock = clock;
  assign brams_4_reset = reset;
  assign brams_4_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_4_io_w_en = io_w_en & io_w_maskOH[4]; // @[SRAM_1.scala 208:37]
  assign brams_4_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_5_clock = clock;
  assign brams_5_reset = reset;
  assign brams_5_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_5_io_w_en = io_w_en & io_w_maskOH[5]; // @[SRAM_1.scala 208:37]
  assign brams_5_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_6_clock = clock;
  assign brams_6_reset = reset;
  assign brams_6_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_6_io_w_en = io_w_en & io_w_maskOH[6]; // @[SRAM_1.scala 208:37]
  assign brams_6_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_7_clock = clock;
  assign brams_7_reset = reset;
  assign brams_7_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_7_io_w_en = io_w_en & io_w_maskOH[7]; // @[SRAM_1.scala 208:37]
  assign brams_7_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  reg  state_8; // @[PRNG.scala 55:49]
  reg  state_9; // @[PRNG.scala 55:49]
  reg  state_10; // @[PRNG.scala 55:49]
  reg  state_11; // @[PRNG.scala 55:49]
  reg  state_12; // @[PRNG.scala 55:49]
  reg  state_13; // @[PRNG.scala 55:49]
  reg  state_14; // @[PRNG.scala 55:49]
  reg  state_15; // @[PRNG.scala 55:49]
  wire  _T_2 = state_15 ^ state_13 ^ state_12 ^ state_10; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  assign io_out_8 = state_8; // @[PRNG.scala 78:10]
  assign io_out_9 = state_9; // @[PRNG.scala 78:10]
  assign io_out_10 = state_10; // @[PRNG.scala 78:10]
  assign io_out_11 = state_11; // @[PRNG.scala 78:10]
  assign io_out_12 = state_12; // @[PRNG.scala 78:10]
  assign io_out_13 = state_13; // @[PRNG.scala 78:10]
  assign io_out_14 = state_14; // @[PRNG.scala 78:10]
  assign io_out_15 = state_15; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T_2; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_4 <= state_3;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_5 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_5 <= state_4;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_6 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_6 <= state_5;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_7 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_7 <= state_6;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_8 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_8 <= state_7;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_9 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_9 <= state_8;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_10 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_10 <= state_9;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_11 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_11 <= state_10;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_12 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_12 <= state_11;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_13 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_13 <= state_12;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_14 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_14 <= state_13;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_15 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_15 <= state_14;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCacheDirectory(
  input         clock,
  input         reset,
  output        io_read_req_ready,
  input         io_read_req_valid,
  input  [31:0] io_read_req_bits_addr,
  output        io_read_resp_bits_hit,
  output [7:0]  io_read_resp_bits_chosenWay,
  output        io_write_req_ready,
  input         io_write_req_valid,
  input  [31:0] io_write_req_bits_addr,
  input  [7:0]  io_write_req_bits_way
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  tagArray_clock; // @[SRAM_1.scala 255:31]
  wire  tagArray_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] tagArray_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  tagArray_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] tagArray_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] tagArray_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  metaArray_clock; // @[SRAM_1.scala 255:31]
  wire  metaArray_reset; // @[SRAM_1.scala 255:31]
  wire [6:0] metaArray_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  metaArray_io_w_en; // @[SRAM_1.scala 255:31]
  wire [6:0] metaArray_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [7:0] metaArray_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  replaceWay_lfsr_prng_clock; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_reset; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_15; // @[PRNG.scala 91:22]
  wire [6:0] rSet = io_read_req_bits_addr[11:5]; // @[Parameters.scala 50:11]
  wire [19:0] rTag = io_read_req_bits_addr[31:12]; // @[Parameters.scala 46:11]
  wire  ren = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  wire [6:0] wSet = io_write_req_bits_addr[11:5]; // @[Parameters.scala 50:11]
  wire [19:0] wTag = io_write_req_bits_addr[31:12]; // @[Parameters.scala 46:11]
  wire  wen = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _T_8 = io_write_req_bits_way[0] + io_write_req_bits_way[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_10 = io_write_req_bits_way[2] + io_write_req_bits_way[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_12 = _T_8 + _T_10; // @[Bitwise.scala 51:90]
  wire [1:0] _T_14 = io_write_req_bits_way[4] + io_write_req_bits_way[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_16 = io_write_req_bits_way[6] + io_write_req_bits_way[7]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_18 = _T_14 + _T_16; // @[Bitwise.scala 51:90]
  wire [3:0] _T_20 = _T_12 + _T_18; // @[Bitwise.scala 51:90]
  wire  _T_46 = ~reset; // @[Directory.scala 69:11]
  wire [19:0] rdata__0 = ren ? tagArray_io_r_data_0 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__1 = ren ? tagArray_io_r_data_1 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__2 = ren ? tagArray_io_r_data_2 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__3 = ren ? tagArray_io_r_data_3 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__4 = ren ? tagArray_io_r_data_4 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__5 = ren ? tagArray_io_r_data_5 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__6 = ren ? tagArray_io_r_data_6 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__7 = ren ? tagArray_io_r_data_7 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_0 = ren ? metaArray_io_r_data_0 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_1 = ren ? metaArray_io_r_data_1 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_2 = ren ? metaArray_io_r_data_2 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_3 = ren ? metaArray_io_r_data_3 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_4 = ren ? metaArray_io_r_data_4 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_5 = ren ? metaArray_io_r_data_5 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_6 = ren ? metaArray_io_r_data_6 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_7 = ren ? metaArray_io_r_data_7 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [15:0] _T_48 = {rdata_1_7,rdata_1_6,rdata_1_5,rdata_1_4,rdata_1_3,rdata_1_2,rdata_1_1,rdata_1_0}; // @[Directory.scala 82:52]
  wire  metaRdVec_0_valid = _T_48[0]; // @[Directory.scala 82:52]
  wire  metaRdVec_1_valid = _T_48[2]; // @[Directory.scala 82:52]
  wire  metaRdVec_2_valid = _T_48[4]; // @[Directory.scala 82:52]
  wire  metaRdVec_3_valid = _T_48[6]; // @[Directory.scala 82:52]
  wire  metaRdVec_4_valid = _T_48[8]; // @[Directory.scala 82:52]
  wire  metaRdVec_5_valid = _T_48[10]; // @[Directory.scala 82:52]
  wire  metaRdVec_6_valid = _T_48[12]; // @[Directory.scala 82:52]
  wire  metaRdVec_7_valid = _T_48[14]; // @[Directory.scala 82:52]
  wire  tagMatchVec_0 = rdata__0 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_1 = rdata__1 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_2 = rdata__2 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_3 = rdata__3 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_4 = rdata__4 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_5 = rdata__5 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_6 = rdata__6 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_7 = rdata__7 == rTag; // @[Directory.scala 85:46]
  wire  _matchWayOH_T = tagMatchVec_0 & metaRdVec_0_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_1 = tagMatchVec_1 & metaRdVec_1_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_2 = tagMatchVec_2 & metaRdVec_2_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_3 = tagMatchVec_3 & metaRdVec_3_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_4 = tagMatchVec_4 & metaRdVec_4_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_5 = tagMatchVec_5 & metaRdVec_5_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_6 = tagMatchVec_6 & metaRdVec_6_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_7 = tagMatchVec_7 & metaRdVec_7_valid; // @[Directory.scala 88:80]
  wire [7:0] matchWayOH = {_matchWayOH_T_7,_matchWayOH_T_6,_matchWayOH_T_5,_matchWayOH_T_4,_matchWayOH_T_3,
    _matchWayOH_T_2,_matchWayOH_T_1,_matchWayOH_T}; // @[Cat.scala 33:92]
  wire  invalidWayVec_0 = ~metaRdVec_0_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_1 = ~metaRdVec_1_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_2 = ~metaRdVec_2_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_3 = ~metaRdVec_3_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_4 = ~metaRdVec_4_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_5 = ~metaRdVec_5_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_6 = ~metaRdVec_6_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_7 = ~metaRdVec_7_valid; // @[Directory.scala 89:53]
  wire [7:0] _invalidWayOH_T_16 = invalidWayVec_6 ? 8'h40 : 8'h80; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_17 = invalidWayVec_5 ? 8'h20 : _invalidWayOH_T_16; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_18 = invalidWayVec_4 ? 8'h10 : _invalidWayOH_T_17; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_19 = invalidWayVec_3 ? 8'h8 : _invalidWayOH_T_18; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_20 = invalidWayVec_2 ? 8'h4 : _invalidWayOH_T_19; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_21 = invalidWayVec_1 ? 8'h2 : _invalidWayOH_T_20; // @[Mux.scala 47:70]
  wire [7:0] invalidWayOH = invalidWayVec_0 ? 8'h1 : _invalidWayOH_T_21; // @[Mux.scala 47:70]
  wire [7:0] _hasInvalidWay_T = {invalidWayVec_0,invalidWayVec_1,invalidWayVec_2,invalidWayVec_3,invalidWayVec_4,
    invalidWayVec_5,invalidWayVec_6,invalidWayVec_7}; // @[Cat.scala 33:92]
  wire  hasInvalidWay = |_hasInvalidWay_T; // @[Directory.scala 91:44]
  wire [7:0] replaceWay_lfsr_lo = {replaceWay_lfsr_prng_io_out_7,replaceWay_lfsr_prng_io_out_6,
    replaceWay_lfsr_prng_io_out_5,replaceWay_lfsr_prng_io_out_4,replaceWay_lfsr_prng_io_out_3,
    replaceWay_lfsr_prng_io_out_2,replaceWay_lfsr_prng_io_out_1,replaceWay_lfsr_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [15:0] replaceWay_lfsr = {replaceWay_lfsr_prng_io_out_15,replaceWay_lfsr_prng_io_out_14,
    replaceWay_lfsr_prng_io_out_13,replaceWay_lfsr_prng_io_out_12,replaceWay_lfsr_prng_io_out_11,
    replaceWay_lfsr_prng_io_out_10,replaceWay_lfsr_prng_io_out_9,replaceWay_lfsr_prng_io_out_8,replaceWay_lfsr_lo}; // @[PRNG.scala 95:17]
  wire [2:0] replaceWay_outputWay_shiftAmount = replaceWay_lfsr[2:0]; // @[DCache.scala 60:39]
  wire [7:0] replaceWay = 8'h1 << replaceWay_outputWay_shiftAmount; // @[OneHot.scala 64:12]
  wire  _replaceWayReg_T = ~io_read_req_valid; // @[Directory.scala 93:65]
  reg [7:0] replaceWayReg; // @[Reg.scala 19:16]
  wire  isHit = |matchWayOH; // @[Directory.scala 95:41]
  wire [7:0] _choseWayOH_T = hasInvalidWay ? invalidWayOH : replaceWayReg; // @[Directory.scala 96:51]
  wire [7:0] choseWayOH = isHit ? matchWayOH : _choseWayOH_T; // @[Directory.scala 96:28]
  wire [1:0] _T_73 = choseWayOH[0] + choseWayOH[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_75 = choseWayOH[2] + choseWayOH[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_77 = _T_73 + _T_75; // @[Bitwise.scala 51:90]
  wire [1:0] _T_79 = choseWayOH[4] + choseWayOH[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_81 = choseWayOH[6] + choseWayOH[7]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_83 = _T_79 + _T_81; // @[Bitwise.scala 51:90]
  wire [3:0] _T_85 = _T_77 + _T_83; // @[Bitwise.scala 51:90]
  SRAMArray_2P_8 tagArray ( // @[SRAM_1.scala 255:31]
    .clock(tagArray_clock),
    .reset(tagArray_reset),
    .io_r_addr(tagArray_io_r_addr),
    .io_r_data_0(tagArray_io_r_data_0),
    .io_r_data_1(tagArray_io_r_data_1),
    .io_r_data_2(tagArray_io_r_data_2),
    .io_r_data_3(tagArray_io_r_data_3),
    .io_r_data_4(tagArray_io_r_data_4),
    .io_r_data_5(tagArray_io_r_data_5),
    .io_r_data_6(tagArray_io_r_data_6),
    .io_r_data_7(tagArray_io_r_data_7),
    .io_w_en(tagArray_io_w_en),
    .io_w_addr(tagArray_io_w_addr),
    .io_w_data_0(tagArray_io_w_data_0),
    .io_w_data_1(tagArray_io_w_data_1),
    .io_w_data_2(tagArray_io_w_data_2),
    .io_w_data_3(tagArray_io_w_data_3),
    .io_w_data_4(tagArray_io_w_data_4),
    .io_w_data_5(tagArray_io_w_data_5),
    .io_w_data_6(tagArray_io_w_data_6),
    .io_w_data_7(tagArray_io_w_data_7),
    .io_w_maskOH(tagArray_io_w_maskOH)
  );
  SRAMArray_2P_9 metaArray ( // @[SRAM_1.scala 255:31]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_addr(metaArray_io_r_addr),
    .io_r_data_0(metaArray_io_r_data_0),
    .io_r_data_1(metaArray_io_r_data_1),
    .io_r_data_2(metaArray_io_r_data_2),
    .io_r_data_3(metaArray_io_r_data_3),
    .io_r_data_4(metaArray_io_r_data_4),
    .io_r_data_5(metaArray_io_r_data_5),
    .io_r_data_6(metaArray_io_r_data_6),
    .io_r_data_7(metaArray_io_r_data_7),
    .io_w_en(metaArray_io_w_en),
    .io_w_addr(metaArray_io_w_addr),
    .io_w_maskOH(metaArray_io_w_maskOH)
  );
  MaxPeriodFibonacciLFSR replaceWay_lfsr_prng ( // @[PRNG.scala 91:22]
    .clock(replaceWay_lfsr_prng_clock),
    .reset(replaceWay_lfsr_prng_reset),
    .io_out_0(replaceWay_lfsr_prng_io_out_0),
    .io_out_1(replaceWay_lfsr_prng_io_out_1),
    .io_out_2(replaceWay_lfsr_prng_io_out_2),
    .io_out_3(replaceWay_lfsr_prng_io_out_3),
    .io_out_4(replaceWay_lfsr_prng_io_out_4),
    .io_out_5(replaceWay_lfsr_prng_io_out_5),
    .io_out_6(replaceWay_lfsr_prng_io_out_6),
    .io_out_7(replaceWay_lfsr_prng_io_out_7),
    .io_out_8(replaceWay_lfsr_prng_io_out_8),
    .io_out_9(replaceWay_lfsr_prng_io_out_9),
    .io_out_10(replaceWay_lfsr_prng_io_out_10),
    .io_out_11(replaceWay_lfsr_prng_io_out_11),
    .io_out_12(replaceWay_lfsr_prng_io_out_12),
    .io_out_13(replaceWay_lfsr_prng_io_out_13),
    .io_out_14(replaceWay_lfsr_prng_io_out_14),
    .io_out_15(replaceWay_lfsr_prng_io_out_15)
  );
  assign io_read_req_ready = 1'h1; // @[Directory.scala 75:29]
  assign io_read_resp_bits_hit = |matchWayOH; // @[Directory.scala 95:41]
  assign io_read_resp_bits_chosenWay = isHit ? matchWayOH : _choseWayOH_T; // @[Directory.scala 96:28]
  assign io_write_req_ready = 1'h1; // @[Directory.scala 76:29]
  assign tagArray_clock = clock;
  assign tagArray_reset = reset;
  assign tagArray_io_r_addr = rSet; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign tagArray_io_w_en = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  assign tagArray_io_w_addr = wSet; // @[Directory.scala 112:15 SRAM_1.scala 237:19]
  assign tagArray_io_w_data_0 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_1 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_2 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_3 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_4 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_5 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_6 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_7 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_maskOH = io_write_req_bits_way; // @[Directory.scala 112:15 SRAM_1.scala 239:21]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r_addr = rSet; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign metaArray_io_w_en = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  assign metaArray_io_w_addr = wSet; // @[Directory.scala 112:15 SRAM_1.scala 237:19]
  assign metaArray_io_w_maskOH = io_write_req_bits_way; // @[Directory.scala 112:15 SRAM_1.scala 239:21]
  assign replaceWay_lfsr_prng_clock = clock;
  assign replaceWay_lfsr_prng_reset = reset;
  always @(posedge clock) begin
    if (_replaceWayReg_T) begin // @[Reg.scala 20:18]
      replaceWayReg <= replaceWay; // @[Reg.scala 20:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_20 < 4'h2)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Error directory write way has multiple valid bit! ==>%d\n    at Directory.scala:69 assert(PopCount(wWay) < 2.U, cf\"Error directory write way has multiple valid bit! ==>${PopCount(wWay)}\")\n"
            ,_T_20); // @[Directory.scala 69:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_20 < 4'h2) & ~reset) begin
          $fatal; // @[Directory.scala 69:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_46 & ~(_T_85 == 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Error chosenWay has multiple valid bit!\n    at Directory.scala:101 assert(PopCount(choseWayOH) === 1.U, \"Error chosenWay has multiple valid bit!\")\n"
            ); // @[Directory.scala 101:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_85 == 4'h1) & _T_46) begin
          $fatal; // @[Directory.scala 101:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wen & _T_46 & ~(_T_20 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: write error, tring to write multiple ways\n    at SRAM_1.scala:235 assert(PopCount(mask) <= 1.U, \"write error, tring to write multiple ways\")\n"
            ); // @[SRAM_1.scala 235:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_20 <= 4'h1) & (wen & _T_46)) begin
          $fatal; // @[SRAM_1.scala 235:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wen & _T_46 & ~(_T_20 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: write error, tring to write multiple ways\n    at SRAM_1.scala:235 assert(PopCount(mask) <= 1.U, \"write error, tring to write multiple ways\")\n"
            ); // @[SRAM_1.scala 235:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_20 <= 4'h1) & (wen & _T_46)) begin
          $fatal; // @[SRAM_1.scala 235:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  replaceWayReg = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RefillPipe(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [31:0]  io_req_bits_addr,
  input  [7:0]   io_req_bits_chosenWay,
  input          io_resp_ready,
  output         io_resp_valid,
  output [31:0]  io_resp_bits_data,
  output [31:0]  io_resp_bits_blockData_0,
  output [31:0]  io_resp_bits_blockData_1,
  output [31:0]  io_resp_bits_blockData_2,
  output [31:0]  io_resp_bits_blockData_3,
  output [31:0]  io_resp_bits_blockData_4,
  output [31:0]  io_resp_bits_blockData_5,
  output [31:0]  io_resp_bits_blockData_6,
  output [31:0]  io_resp_bits_blockData_7,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [127:0] io_tlbus_req_bits_size,
  output [31:0]  io_tlbus_req_bits_address,
  output         io_tlbus_resp_ready,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data,
  output         io_dirWrite_req_valid,
  output [31:0]  io_dirWrite_req_bits_addr,
  output [7:0]   io_dirWrite_req_bits_way,
  output         io_dataWrite_req_valid,
  output [6:0]   io_dataWrite_req_bits_set,
  output [31:0]  io_dataWrite_req_bits_data_0,
  output [31:0]  io_dataWrite_req_bits_data_1,
  output [31:0]  io_dataWrite_req_bits_data_2,
  output [31:0]  io_dataWrite_req_bits_data_3,
  output [31:0]  io_dataWrite_req_bits_data_4,
  output [31:0]  io_dataWrite_req_bits_data_5,
  output [31:0]  io_dataWrite_req_bits_data_6,
  output [31:0]  io_dataWrite_req_bits_data_7,
  output [7:0]   io_dataWrite_req_bits_blockMask,
  output [7:0]   io_dataWrite_req_bits_way
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[RefillPipe.scala 42:24]
  wire  _io_req_ready_T = state == 2'h0; // @[RefillPipe.scala 45:27]
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] reqReg_addr; // @[Reg.scala 19:16]
  reg [7:0] reqReg_chosenWay; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  reg  reqValidReg; // @[Reg.scala 19:16]
  wire  _GEN_2 = _reqReg_T | reqValidReg; // @[Reg.scala 19:16 20:{18,22}]
  wire [7:0] dataBlockSelOH = 8'h1 << reqReg_addr[4:2]; // @[OneHot.scala 57:35]
  reg  beatCounter_value; // @[Counter.scala 61:40]
  wire [1:0] beatOH = 2'h1 << beatCounter_value; // @[OneHot.scala 64:12]
  wire  _refillFire_T = io_tlbus_resp_ready & io_tlbus_resp_valid; // @[Decoupled.scala 51:35]
  wire  refillFire = _refillFire_T & io_tlbus_resp_bits_opcode == 3'h1; // @[RefillPipe.scala 59:41]
  wire  refillLastBeat = refillFire & beatCounter_value; // @[RefillPipe.scala 60:37]
  wire  _T_2 = io_tlbus_req_ready & io_tlbus_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_4 = _T_2 ? 2'h2 : {{1'd0}, _reqReg_T}; // @[RefillPipe.scala 71:33 72:23]
  wire  _GEN_5 = _T_2 ? 1'h0 : _GEN_2; // @[RefillPipe.scala 71:33 73:25]
  wire [1:0] _GEN_6 = _io_req_ready_T ? _GEN_4 : 2'h0; // @[RefillPipe.scala 66:27 43:29]
  wire  _GEN_7 = _io_req_ready_T ? _GEN_5 : _GEN_2; // @[RefillPipe.scala 66:27]
  wire [1:0] _GEN_8 = _T_2 ? 2'h2 : 2'h1; // @[RefillPipe.scala 80:19 81:33 82:23]
  wire  _T_5 = state == 2'h2; // @[RefillPipe.scala 89:16]
  wire [1:0] _GEN_12 = io_resp_valid ? 2'h0 : 2'h3; // @[RefillPipe.scala 92:23 93:32 94:27]
  wire  _T_7 = state == 2'h3; // @[RefillPipe.scala 105:16]
  wire  refillSafe = refillFire & _T_5; // @[RefillPipe.scala 115:33]
  wire [3:0] _blockMask_T_3 = beatOH[0] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _blockMask_T_5 = beatOH[1] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [255:0] _T_9 = {io_tlbus_resp_bits_data,io_tlbus_resp_bits_data}; // @[Cat.scala 33:92]
  reg [31:0] refillBlockDataArray_0_0; // @[RefillPipe.scala 133:39]
  reg [31:0] refillBlockDataArray_0_1; // @[RefillPipe.scala 133:39]
  reg [31:0] refillBlockDataArray_0_2; // @[RefillPipe.scala 133:39]
  reg [31:0] refillBlockDataArray_0_3; // @[RefillPipe.scala 133:39]
  wire [255:0] _io_resp_bits_data_T = {io_tlbus_resp_bits_data,refillBlockDataArray_0_3,refillBlockDataArray_0_2,
    refillBlockDataArray_0_1,refillBlockDataArray_0_0}; // @[RefillPipe.scala 141:72]
  wire [31:0] _io_resp_bits_data_T_17 = dataBlockSelOH[0] ? _io_resp_bits_data_T[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_18 = dataBlockSelOH[1] ? _io_resp_bits_data_T[63:32] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_19 = dataBlockSelOH[2] ? _io_resp_bits_data_T[95:64] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_20 = dataBlockSelOH[3] ? _io_resp_bits_data_T[127:96] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_21 = dataBlockSelOH[4] ? _io_resp_bits_data_T[159:128] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_22 = dataBlockSelOH[5] ? _io_resp_bits_data_T[191:160] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_23 = dataBlockSelOH[6] ? _io_resp_bits_data_T[223:192] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_24 = dataBlockSelOH[7] ? _io_resp_bits_data_T[255:224] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_25 = _io_resp_bits_data_T_17 | _io_resp_bits_data_T_18; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_26 = _io_resp_bits_data_T_25 | _io_resp_bits_data_T_19; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_27 = _io_resp_bits_data_T_26 | _io_resp_bits_data_T_20; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_28 = _io_resp_bits_data_T_27 | _io_resp_bits_data_T_21; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_29 = _io_resp_bits_data_T_28 | _io_resp_bits_data_T_22; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_30 = _io_resp_bits_data_T_29 | _io_resp_bits_data_T_23; // @[Mux.scala 27:73]
  reg [63:0] c; // @[util.scala 162:24]
  wire [63:0] _c_T_1 = c + 64'h1; // @[util.scala 163:16]
  reg [63:0] c_1; // @[util.scala 162:24]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[util.scala 163:16]
  assign io_req_ready = state == 2'h0; // @[RefillPipe.scala 45:27]
  assign io_resp_valid = _T_7 | refillLastBeat; // @[RefillPipe.scala 140:38]
  assign io_resp_bits_data = _io_resp_bits_data_T_30 | _io_resp_bits_data_T_24; // @[Mux.scala 27:73]
  assign io_resp_bits_blockData_0 = _io_resp_bits_data_T[31:0]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_1 = _io_resp_bits_data_T[63:32]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_2 = _io_resp_bits_data_T[95:64]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_3 = _io_resp_bits_data_T[127:96]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_4 = _io_resp_bits_data_T[159:128]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_5 = _io_resp_bits_data_T[191:160]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_6 = _io_resp_bits_data_T[223:192]; // @[RefillPipe.scala 142:55]
  assign io_resp_bits_blockData_7 = _io_resp_bits_data_T[255:224]; // @[RefillPipe.scala 142:55]
  assign io_tlbus_req_valid = _reqReg_T | reqValidReg; // @[RefillPipe.scala 50:23]
  assign io_tlbus_req_bits_size = 128'h20; // @[RefillPipe.scala 150:28]
  assign io_tlbus_req_bits_address = {_GEN_0[31:5],5'h0}; // @[Cat.scala 33:92]
  assign io_tlbus_resp_ready = 1'h1; // @[RefillPipe.scala 62:51]
  assign io_dirWrite_req_valid = refillSafe & beatCounter_value; // @[RefillPipe.scala 116:41]
  assign io_dirWrite_req_bits_addr = reqReg_addr; // @[RefillPipe.scala 117:31]
  assign io_dirWrite_req_bits_way = reqReg_chosenWay; // @[RefillPipe.scala 122:30]
  assign io_dataWrite_req_valid = refillFire & _T_5; // @[RefillPipe.scala 115:33]
  assign io_dataWrite_req_bits_set = reqReg_addr[11:5]; // @[Parameters.scala 50:11]
  assign io_dataWrite_req_bits_data_0 = _T_9[31:0]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_1 = _T_9[63:32]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_2 = _T_9[95:64]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_3 = _T_9[127:96]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_4 = _T_9[159:128]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_5 = _T_9[191:160]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_6 = _T_9[223:192]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_7 = _T_9[255:224]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_blockMask = {_blockMask_T_5,_blockMask_T_3}; // @[Cat.scala 33:92]
  assign io_dataWrite_req_bits_way = reqReg_chosenWay; // @[RefillPipe.scala 128:31]
  always @(posedge clock) begin
    if (reset) begin // @[RefillPipe.scala 42:24]
      state <= 2'h0; // @[RefillPipe.scala 42:24]
    end else if (state == 2'h3) begin // @[RefillPipe.scala 105:27]
      state <= _GEN_12;
    end else if (state == 2'h2) begin // @[RefillPipe.scala 89:33]
      if (refillLastBeat) begin // @[RefillPipe.scala 91:30]
        state <= _GEN_12;
      end else begin
        state <= 2'h2;
      end
    end else if (state == 2'h1) begin // @[RefillPipe.scala 79:26]
      state <= _GEN_8;
    end else begin
      state <= _GEN_6;
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_addr <= io_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_chosenWay <= io_req_bits_chosenWay; // @[Reg.scala 20:22]
    end
    if (state == 2'h1) begin // @[RefillPipe.scala 79:26]
      if (_T_2) begin // @[RefillPipe.scala 81:33]
        reqValidReg <= 1'h0; // @[RefillPipe.scala 83:25]
      end else begin
        reqValidReg <= _GEN_7;
      end
    end else begin
      reqValidReg <= _GEN_7;
    end
    if (reset) begin // @[Counter.scala 61:40]
      beatCounter_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (state == 2'h2) begin // @[RefillPipe.scala 89:33]
      if (refillLastBeat) begin // @[RefillPipe.scala 91:30]
        beatCounter_value <= 1'h0; // @[Counter.scala 98:11]
      end else if (refillFire) begin // @[RefillPipe.scala 97:32]
        beatCounter_value <= beatCounter_value + 1'h1; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[RefillPipe.scala 133:39]
      refillBlockDataArray_0_0 <= 32'h0; // @[RefillPipe.scala 133:39]
    end else if (refillFire) begin // @[RefillPipe.scala 134:22]
      if (~beatCounter_value) begin // @[RefillPipe.scala 135:49]
        refillBlockDataArray_0_0 <= io_tlbus_resp_bits_data[31:0]; // @[RefillPipe.scala 135:49]
      end
    end
    if (reset) begin // @[RefillPipe.scala 133:39]
      refillBlockDataArray_0_1 <= 32'h0; // @[RefillPipe.scala 133:39]
    end else if (refillFire) begin // @[RefillPipe.scala 134:22]
      if (~beatCounter_value) begin // @[RefillPipe.scala 135:49]
        refillBlockDataArray_0_1 <= io_tlbus_resp_bits_data[63:32]; // @[RefillPipe.scala 135:49]
      end
    end
    if (reset) begin // @[RefillPipe.scala 133:39]
      refillBlockDataArray_0_2 <= 32'h0; // @[RefillPipe.scala 133:39]
    end else if (refillFire) begin // @[RefillPipe.scala 134:22]
      if (~beatCounter_value) begin // @[RefillPipe.scala 135:49]
        refillBlockDataArray_0_2 <= io_tlbus_resp_bits_data[95:64]; // @[RefillPipe.scala 135:49]
      end
    end
    if (reset) begin // @[RefillPipe.scala 133:39]
      refillBlockDataArray_0_3 <= 32'h0; // @[RefillPipe.scala 133:39]
    end else if (refillFire) begin // @[RefillPipe.scala 134:22]
      if (~beatCounter_value) begin // @[RefillPipe.scala 135:49]
        refillBlockDataArray_0_3 <= io_tlbus_resp_bits_data[127:96]; // @[RefillPipe.scala 135:49]
      end
    end
    if (reset) begin // @[util.scala 162:24]
      c <= 64'h0; // @[util.scala 162:24]
    end else begin
      c <= _c_T_1; // @[util.scala 163:11]
    end
    if (reset) begin // @[util.scala 162:24]
      c_1 <= 64'h0; // @[util.scala 162:24]
    end else begin
      c_1 <= _c_T_3; // @[util.scala 163:11]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [RefillPipe] req ==> addr: 0x%x size:%d\n",c,
            io_tlbus_req_bits_address,io_tlbus_req_bits_size); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (refillFire & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [RefillPipe] resp <== data: 0x%x beat: %d\n",c_1,
            io_tlbus_resp_bits_data,beatCounter_value); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reqReg_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqReg_chosenWay = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  reqValidReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  beatCounter_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  refillBlockDataArray_0_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  refillBlockDataArray_0_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  refillBlockDataArray_0_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  refillBlockDataArray_0_3 = _RAND_8[31:0];
  _RAND_9 = {2{`RANDOM}};
  c = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  c_1 = _RAND_10[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RefillBuffer(
  input          clock,
  input          reset,
  input          io_write_valid,
  input  [31:0]  io_write_bits_cacheLineAddr,
  input  [127:0] io_write_bits_data,
  output [31:0]  io_read_cacheLineAddr_0,
  output [31:0]  io_read_cacheLineAddr_1,
  output [31:0]  io_read_cacheLineData_0_0,
  output [31:0]  io_read_cacheLineData_0_1,
  output [31:0]  io_read_cacheLineData_0_2,
  output [31:0]  io_read_cacheLineData_0_3,
  output [31:0]  io_read_cacheLineData_0_4,
  output [31:0]  io_read_cacheLineData_0_5,
  output [31:0]  io_read_cacheLineData_0_6,
  output [31:0]  io_read_cacheLineData_0_7,
  output [31:0]  io_read_cacheLineData_1_0,
  output [31:0]  io_read_cacheLineData_1_1,
  output [31:0]  io_read_cacheLineData_1_2,
  output [31:0]  io_read_cacheLineData_1_3,
  output [31:0]  io_read_cacheLineData_1_4,
  output [31:0]  io_read_cacheLineData_1_5,
  output [31:0]  io_read_cacheLineData_1_6,
  output [31:0]  io_read_cacheLineData_1_7,
  output         io_read_valids_0,
  output         io_read_valids_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] buf_0_0; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_1; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_2; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_3; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_4; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_5; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_6; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_0_7; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_0; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_1; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_2; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_3; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_4; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_5; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_6; // @[RefillBuffer.scala 23:18]
  reg [31:0] buf_1_7; // @[RefillBuffer.scala 23:18]
  reg [31:0] addr_0; // @[RefillBuffer.scala 24:19]
  reg [31:0] addr_1; // @[RefillBuffer.scala 24:19]
  reg  wrPtr_value; // @[Counter.scala 61:40]
  reg  beatCounter_value; // @[Counter.scala 61:40]
  wire [31:0] _addr_T_2 = {io_write_bits_cacheLineAddr[31:5],5'h0}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_60 = {{1'd0}, beatCounter_value}; // @[RefillBuffer.scala 23:18 43:{45,45}]
  wire [2:0] _GEN_66 = {{2'd0}, beatCounter_value}; // @[RefillBuffer.scala 23:18 43:{45,45}]
  assign io_read_cacheLineAddr_0 = addr_0; // @[RefillBuffer.scala 47:27]
  assign io_read_cacheLineAddr_1 = addr_1; // @[RefillBuffer.scala 47:27]
  assign io_read_cacheLineData_0_0 = buf_0_0; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_1 = buf_0_1; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_2 = buf_0_2; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_3 = buf_0_3; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_4 = buf_0_4; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_5 = buf_0_5; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_6 = buf_0_6; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_0_7 = buf_0_7; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_0 = buf_1_0; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_1 = buf_1_1; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_2 = buf_1_2; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_3 = buf_1_3; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_4 = buf_1_4; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_5 = buf_1_5; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_6 = buf_1_6; // @[RefillBuffer.scala 48:27]
  assign io_read_cacheLineData_1_7 = buf_1_7; // @[RefillBuffer.scala 48:27]
  assign io_read_valids_0 = 1'h0; // @[RefillBuffer.scala 49:20]
  assign io_read_valids_1 = 1'h0; // @[RefillBuffer.scala 49:20]
  always @(posedge clock) begin
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & ~beatCounter_value) begin // @[RefillBuffer.scala 43:45]
        buf_0_0 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & beatCounter_value) begin // @[RefillBuffer.scala 43:45]
        buf_0_1 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 2'h2 == _GEN_60) begin // @[RefillBuffer.scala 43:45]
        buf_0_2 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 2'h3 == _GEN_60) begin // @[RefillBuffer.scala 43:45]
        buf_0_3 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 3'h4 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_0_4 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 3'h5 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_0_5 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 3'h6 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_0_6 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (~wrPtr_value & 3'h7 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_0_7 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & ~beatCounter_value) begin // @[RefillBuffer.scala 43:45]
        buf_1_0 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & beatCounter_value) begin // @[RefillBuffer.scala 43:45]
        buf_1_1 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 2'h2 == _GEN_60) begin // @[RefillBuffer.scala 43:45]
        buf_1_2 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 2'h3 == _GEN_60) begin // @[RefillBuffer.scala 43:45]
        buf_1_3 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 3'h4 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_1_4 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 3'h5 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_1_5 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 3'h6 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_1_6 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid) begin // @[RefillBuffer.scala 42:25]
      if (wrPtr_value & 3'h7 == _GEN_66) begin // @[RefillBuffer.scala 43:45]
        buf_1_7 <= io_write_bits_data[31:0]; // @[RefillBuffer.scala 43:45]
      end
    end
    if (io_write_valid & beatCounter_value) begin // @[RefillBuffer.scala 34:37]
      if (~wrPtr_value) begin // @[RefillBuffer.scala 37:27]
        addr_0 <= _addr_T_2; // @[RefillBuffer.scala 37:27]
      end
    end
    if (io_write_valid & beatCounter_value) begin // @[RefillBuffer.scala 34:37]
      if (wrPtr_value) begin // @[RefillBuffer.scala 37:27]
        addr_1 <= _addr_T_2; // @[RefillBuffer.scala 37:27]
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      wrPtr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (io_write_valid & beatCounter_value) begin // @[RefillBuffer.scala 34:37]
      wrPtr_value <= wrPtr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      beatCounter_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (io_write_valid & beatCounter_value) begin // @[RefillBuffer.scala 34:37]
      beatCounter_value <= 1'h0; // @[Counter.scala 98:11]
    end else if (io_write_valid) begin // @[RefillBuffer.scala 38:31]
      beatCounter_value <= beatCounter_value + 1'h1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buf_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  buf_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  buf_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  buf_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  buf_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  buf_0_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  buf_0_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  buf_0_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  buf_1_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  buf_1_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  buf_1_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  buf_1_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  buf_1_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  buf_1_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  buf_1_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  buf_1_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  addr_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  addr_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  wrPtr_value = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  beatCounter_value = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input          clock,
  input          reset,
  output         io_read_req_ready,
  input          io_read_req_valid,
  input  [31:0]  io_read_req_bits_addr,
  input          io_read_resp_ready,
  output         io_read_resp_valid,
  output [31:0]  io_read_resp_bits_data,
  output [31:0]  io_read_resp_bits_inst_0,
  output [31:0]  io_read_resp_bits_inst_1,
  output [31:0]  io_read_resp_bits_inst_2,
  output [31:0]  io_read_resp_bits_inst_3,
  output [2:0]   io_read_resp_bits_size,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [31:0]  io_tlbus_req_bits_address,
  output         io_tlbus_resp_ready,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
`endif // RANDOMIZE_REG_INIT
  wire  db_clock; // @[ICache.scala 56:20]
  wire  db_reset; // @[ICache.scala 56:20]
  wire  db_io_read_req_ready; // @[ICache.scala 56:20]
  wire  db_io_read_req_valid; // @[ICache.scala 56:20]
  wire [6:0] db_io_read_req_bits_set; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_0_0; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_0_1; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_0_2; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_0_3; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_0_4; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_0_5; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_0_6; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_0_7; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_1_0; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_1_1; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_1_2; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_1_3; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_1_4; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_1_5; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_1_6; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_1_7; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_2_0; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_2_1; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_2_2; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_2_3; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_2_4; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_2_5; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_2_6; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_2_7; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_3_0; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_3_1; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_3_2; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_3_3; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_3_4; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_3_5; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_3_6; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_3_7; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_4_0; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_4_1; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_4_2; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_4_3; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_4_4; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_4_5; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_4_6; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_4_7; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_5_0; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_5_1; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_5_2; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_5_3; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_5_4; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_5_5; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_5_6; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_5_7; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_6_0; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_6_1; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_6_2; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_6_3; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_6_4; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_6_5; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_6_6; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_6_7; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_7_0; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_7_1; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_7_2; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_7_3; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_7_4; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_7_5; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_7_6; // @[ICache.scala 56:20]
  wire [31:0] db_io_read_resp_7_7; // @[ICache.scala 56:20]
  wire  db_io_write_req_ready; // @[ICache.scala 56:20]
  wire  db_io_write_req_valid; // @[ICache.scala 56:20]
  wire [6:0] db_io_write_req_bits_set; // @[ICache.scala 56:20]
  wire [31:0] db_io_write_req_bits_data_0; // @[ICache.scala 56:20]
  wire [31:0] db_io_write_req_bits_data_1; // @[ICache.scala 56:20]
  wire [31:0] db_io_write_req_bits_data_2; // @[ICache.scala 56:20]
  wire [31:0] db_io_write_req_bits_data_3; // @[ICache.scala 56:20]
  wire [31:0] db_io_write_req_bits_data_4; // @[ICache.scala 56:20]
  wire [31:0] db_io_write_req_bits_data_5; // @[ICache.scala 56:20]
  wire [31:0] db_io_write_req_bits_data_6; // @[ICache.scala 56:20]
  wire [31:0] db_io_write_req_bits_data_7; // @[ICache.scala 56:20]
  wire [7:0] db_io_write_req_bits_blockMask; // @[ICache.scala 56:20]
  wire [7:0] db_io_write_req_bits_way; // @[ICache.scala 56:20]
  wire  dir_clock; // @[ICache.scala 57:21]
  wire  dir_reset; // @[ICache.scala 57:21]
  wire  dir_io_read_req_ready; // @[ICache.scala 57:21]
  wire  dir_io_read_req_valid; // @[ICache.scala 57:21]
  wire [31:0] dir_io_read_req_bits_addr; // @[ICache.scala 57:21]
  wire  dir_io_read_resp_bits_hit; // @[ICache.scala 57:21]
  wire [7:0] dir_io_read_resp_bits_chosenWay; // @[ICache.scala 57:21]
  wire  dir_io_write_req_ready; // @[ICache.scala 57:21]
  wire  dir_io_write_req_valid; // @[ICache.scala 57:21]
  wire [31:0] dir_io_write_req_bits_addr; // @[ICache.scala 57:21]
  wire [7:0] dir_io_write_req_bits_way; // @[ICache.scala 57:21]
  wire  refillPipe_clock; // @[ICache.scala 58:28]
  wire  refillPipe_reset; // @[ICache.scala 58:28]
  wire  refillPipe_io_req_ready; // @[ICache.scala 58:28]
  wire  refillPipe_io_req_valid; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_req_bits_addr; // @[ICache.scala 58:28]
  wire [7:0] refillPipe_io_req_bits_chosenWay; // @[ICache.scala 58:28]
  wire  refillPipe_io_resp_ready; // @[ICache.scala 58:28]
  wire  refillPipe_io_resp_valid; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_resp_bits_data; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_0; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_1; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_2; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_3; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_4; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_5; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_6; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_resp_bits_blockData_7; // @[ICache.scala 58:28]
  wire  refillPipe_io_tlbus_req_ready; // @[ICache.scala 58:28]
  wire  refillPipe_io_tlbus_req_valid; // @[ICache.scala 58:28]
  wire [127:0] refillPipe_io_tlbus_req_bits_size; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_tlbus_req_bits_address; // @[ICache.scala 58:28]
  wire  refillPipe_io_tlbus_resp_ready; // @[ICache.scala 58:28]
  wire  refillPipe_io_tlbus_resp_valid; // @[ICache.scala 58:28]
  wire [2:0] refillPipe_io_tlbus_resp_bits_opcode; // @[ICache.scala 58:28]
  wire [127:0] refillPipe_io_tlbus_resp_bits_data; // @[ICache.scala 58:28]
  wire  refillPipe_io_dirWrite_req_valid; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_dirWrite_req_bits_addr; // @[ICache.scala 58:28]
  wire [7:0] refillPipe_io_dirWrite_req_bits_way; // @[ICache.scala 58:28]
  wire  refillPipe_io_dataWrite_req_valid; // @[ICache.scala 58:28]
  wire [6:0] refillPipe_io_dataWrite_req_bits_set; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_0; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_1; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_2; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_3; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_4; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_5; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_6; // @[ICache.scala 58:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_7; // @[ICache.scala 58:28]
  wire [7:0] refillPipe_io_dataWrite_req_bits_blockMask; // @[ICache.scala 58:28]
  wire [7:0] refillPipe_io_dataWrite_req_bits_way; // @[ICache.scala 58:28]
  wire  refillBuffer_clock; // @[ICache.scala 65:30]
  wire  refillBuffer_reset; // @[ICache.scala 65:30]
  wire  refillBuffer_io_write_valid; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_write_bits_cacheLineAddr; // @[ICache.scala 65:30]
  wire [127:0] refillBuffer_io_write_bits_data; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineAddr_0; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineAddr_1; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_0; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_1; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_2; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_3; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_4; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_5; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_6; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_0_7; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_0; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_1; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_2; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_3; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_4; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_5; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_6; // @[ICache.scala 65:30]
  wire [31:0] refillBuffer_io_read_cacheLineData_1_7; // @[ICache.scala 65:30]
  wire  refillBuffer_io_read_valids_0; // @[ICache.scala 65:30]
  wire  refillBuffer_io_read_valids_1; // @[ICache.scala 65:30]
  reg  s0_full; // @[ICache.scala 75:26]
  wire  s0_latch = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  reg  s1_full; // @[ICache.scala 112:26]
  reg  s1_info_dirInfo_hit; // @[Reg.scala 19:16]
  wire  _s1_valid_T_2 = ~s1_info_dirInfo_hit; // @[ICache.scala 137:25]
  wire  _s1_valid_T_3 = refillPipe_io_req_ready & refillPipe_io_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] s1_info_req_addr; // @[Reg.scala 19:16]
  wire [31:0] _bypassVec_T_2 = {s1_info_req_addr[31:5],5'h0}; // @[Cat.scala 33:92]
  wire  bypassVec_0 = refillBuffer_io_read_cacheLineAddr_0 == _bypassVec_T_2 & refillBuffer_io_read_valids_0; // @[ICache.scala 124:154]
  wire  bypassVec_1 = refillBuffer_io_read_cacheLineAddr_1 == _bypassVec_T_2 & refillBuffer_io_read_valids_1; // @[ICache.scala 124:154]
  wire [1:0] _s1_bypass_T = {bypassVec_0,bypassVec_1}; // @[Cat.scala 33:92]
  wire  s1_bypass = |_s1_bypass_T & s1_full & _s1_valid_T_2; // @[ICache.scala 125:51]
  wire  _s1_valid_T_5 = ~s1_bypass; // @[ICache.scala 137:75]
  wire  _s1_valid_T_6 = ~s1_info_dirInfo_hit & _s1_valid_T_3 & ~s1_bypass; // @[ICache.scala 137:72]
  wire  _s1_valid_T_7 = s1_info_dirInfo_hit & io_read_resp_valid | _s1_valid_T_6; // @[ICache.scala 136:71]
  wire  _s1_valid_T_11 = _s1_valid_T_2 & s1_bypass & io_read_resp_valid; // @[ICache.scala 138:59]
  wire  _s1_valid_T_12 = _s1_valid_T_7 | _s1_valid_T_11; // @[ICache.scala 137:86]
  wire  s1_valid = s1_full & _s1_valid_T_12; // @[ICache.scala 136:25]
  reg  s2_full; // @[ICache.scala 144:26]
  reg  s2_dirInfo_hit; // @[Reg.scala 19:16]
  wire  _s2_valid_T = ~s2_dirInfo_hit; // @[ICache.scala 163:47]
  reg  s2_bypass; // @[Reg.scala 19:16]
  wire  s2_fire = s2_full & (s2_dirInfo_hit | ~s2_dirInfo_hit & io_read_resp_valid | s2_bypass); // @[ICache.scala 163:25]
  wire  s2_ready = ~s2_full | s2_fire; // @[ICache.scala 150:26]
  wire  s1_fire = s1_valid & s2_ready; // @[ICache.scala 114:28]
  wire  s1_ready = ~s1_full | s1_fire; // @[ICache.scala 119:26]
  wire  s0_fire = s0_full & s1_ready; // @[ICache.scala 77:28]
  reg [31:0] s0_req_r_addr; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = s0_latch ? io_read_req_bits_addr : s0_req_r_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_1 = s0_full & s0_fire ? 1'h0 : s0_full; // @[ICache.scala 75:26 83:{35,45}]
  wire  _GEN_2 = s0_latch | _GEN_1; // @[ICache.scala 82:{20,30}]
  reg [7:0] s1_info_dirInfo_chosenWay; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_0_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_1_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_2_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_3_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_4_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_5_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_6_7; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_0; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_1; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_2; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_3; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_4; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_5; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_6; // @[Reg.scala 19:16]
  reg [31:0] s1_info_rdData_7_7; // @[Reg.scala 19:16]
  wire [31:0] s0_info_rdData_0_0 = db_io_read_resp_0_0; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_0_1 = db_io_read_resp_0_1; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_0_2 = db_io_read_resp_0_2; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_0_3 = db_io_read_resp_0_3; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_0_4 = db_io_read_resp_0_4; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_0_5 = db_io_read_resp_0_5; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_0_6 = db_io_read_resp_0_6; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_0_7 = db_io_read_resp_0_7; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_1_0 = db_io_read_resp_1_0; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_1_1 = db_io_read_resp_1_1; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_1_2 = db_io_read_resp_1_2; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_1_3 = db_io_read_resp_1_3; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_1_4 = db_io_read_resp_1_4; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_1_5 = db_io_read_resp_1_5; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_1_6 = db_io_read_resp_1_6; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_1_7 = db_io_read_resp_1_7; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_2_0 = db_io_read_resp_2_0; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_2_1 = db_io_read_resp_2_1; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_2_2 = db_io_read_resp_2_2; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_2_3 = db_io_read_resp_2_3; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_2_4 = db_io_read_resp_2_4; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_2_5 = db_io_read_resp_2_5; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_2_6 = db_io_read_resp_2_6; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_2_7 = db_io_read_resp_2_7; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_3_0 = db_io_read_resp_3_0; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_3_1 = db_io_read_resp_3_1; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_3_2 = db_io_read_resp_3_2; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_3_3 = db_io_read_resp_3_3; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_3_4 = db_io_read_resp_3_4; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_3_5 = db_io_read_resp_3_5; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_3_6 = db_io_read_resp_3_6; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_3_7 = db_io_read_resp_3_7; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_4_0 = db_io_read_resp_4_0; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_4_1 = db_io_read_resp_4_1; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_4_2 = db_io_read_resp_4_2; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_4_3 = db_io_read_resp_4_3; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_4_4 = db_io_read_resp_4_4; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_4_5 = db_io_read_resp_4_5; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_4_6 = db_io_read_resp_4_6; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_4_7 = db_io_read_resp_4_7; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_5_0 = db_io_read_resp_5_0; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_5_1 = db_io_read_resp_5_1; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_5_2 = db_io_read_resp_5_2; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_5_3 = db_io_read_resp_5_3; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_5_4 = db_io_read_resp_5_4; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_5_5 = db_io_read_resp_5_5; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_5_6 = db_io_read_resp_5_6; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_5_7 = db_io_read_resp_5_7; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_6_0 = db_io_read_resp_6_0; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_6_1 = db_io_read_resp_6_1; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_6_2 = db_io_read_resp_6_2; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_6_3 = db_io_read_resp_6_3; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_6_4 = db_io_read_resp_6_4; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_6_5 = db_io_read_resp_6_5; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_6_6 = db_io_read_resp_6_6; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_6_7 = db_io_read_resp_6_7; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_7_0 = db_io_read_resp_7_0; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_7_1 = db_io_read_resp_7_1; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_7_2 = db_io_read_resp_7_2; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_7_3 = db_io_read_resp_7_3; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_7_4 = db_io_read_resp_7_4; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_7_5 = db_io_read_resp_7_5; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_7_6 = db_io_read_resp_7_6; // @[ICache.scala 103:23 106:20]
  wire [31:0] s0_info_rdData_7_7 = db_io_read_resp_7_7; // @[ICache.scala 103:23 106:20]
  wire  s0_info_dirInfo_hit = dir_io_read_resp_bits_hit; // @[ICache.scala 103:23 104:21]
  wire [7:0] s0_info_dirInfo_chosenWay = dir_io_read_resp_bits_chosenWay; // @[ICache.scala 103:23 104:21]
  wire [7:0] s1_blockSel = 8'h1 << s1_info_req_addr[4:2]; // @[OneHot.scala 57:35]
  wire [31:0] _s1_rdBlockData_T_8 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_9 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_10 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_11 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_12 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_13 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_14 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_15 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_16 = _s1_rdBlockData_T_8 | _s1_rdBlockData_T_9; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_17 = _s1_rdBlockData_T_16 | _s1_rdBlockData_T_10; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_18 = _s1_rdBlockData_T_17 | _s1_rdBlockData_T_11; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_19 = _s1_rdBlockData_T_18 | _s1_rdBlockData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_20 = _s1_rdBlockData_T_19 | _s1_rdBlockData_T_13; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_21 = _s1_rdBlockData_T_20 | _s1_rdBlockData_T_14; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_0 = _s1_rdBlockData_T_21 | _s1_rdBlockData_T_15; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_23 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_24 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_25 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_26 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_27 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_28 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_29 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_30 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_31 = _s1_rdBlockData_T_23 | _s1_rdBlockData_T_24; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_32 = _s1_rdBlockData_T_31 | _s1_rdBlockData_T_25; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_33 = _s1_rdBlockData_T_32 | _s1_rdBlockData_T_26; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_34 = _s1_rdBlockData_T_33 | _s1_rdBlockData_T_27; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_35 = _s1_rdBlockData_T_34 | _s1_rdBlockData_T_28; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_36 = _s1_rdBlockData_T_35 | _s1_rdBlockData_T_29; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_1 = _s1_rdBlockData_T_36 | _s1_rdBlockData_T_30; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_38 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_39 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_40 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_41 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_42 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_43 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_44 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_45 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_46 = _s1_rdBlockData_T_38 | _s1_rdBlockData_T_39; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_47 = _s1_rdBlockData_T_46 | _s1_rdBlockData_T_40; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_48 = _s1_rdBlockData_T_47 | _s1_rdBlockData_T_41; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_49 = _s1_rdBlockData_T_48 | _s1_rdBlockData_T_42; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_50 = _s1_rdBlockData_T_49 | _s1_rdBlockData_T_43; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_51 = _s1_rdBlockData_T_50 | _s1_rdBlockData_T_44; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_2 = _s1_rdBlockData_T_51 | _s1_rdBlockData_T_45; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_53 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_54 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_55 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_56 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_57 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_58 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_59 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_60 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_61 = _s1_rdBlockData_T_53 | _s1_rdBlockData_T_54; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_62 = _s1_rdBlockData_T_61 | _s1_rdBlockData_T_55; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_63 = _s1_rdBlockData_T_62 | _s1_rdBlockData_T_56; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_64 = _s1_rdBlockData_T_63 | _s1_rdBlockData_T_57; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_65 = _s1_rdBlockData_T_64 | _s1_rdBlockData_T_58; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_66 = _s1_rdBlockData_T_65 | _s1_rdBlockData_T_59; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_3 = _s1_rdBlockData_T_66 | _s1_rdBlockData_T_60; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_68 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_69 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_70 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_71 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_72 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_73 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_74 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_75 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_76 = _s1_rdBlockData_T_68 | _s1_rdBlockData_T_69; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_77 = _s1_rdBlockData_T_76 | _s1_rdBlockData_T_70; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_78 = _s1_rdBlockData_T_77 | _s1_rdBlockData_T_71; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_79 = _s1_rdBlockData_T_78 | _s1_rdBlockData_T_72; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_80 = _s1_rdBlockData_T_79 | _s1_rdBlockData_T_73; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_81 = _s1_rdBlockData_T_80 | _s1_rdBlockData_T_74; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_4 = _s1_rdBlockData_T_81 | _s1_rdBlockData_T_75; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_83 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_84 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_85 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_86 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_87 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_88 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_89 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_90 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_91 = _s1_rdBlockData_T_83 | _s1_rdBlockData_T_84; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_92 = _s1_rdBlockData_T_91 | _s1_rdBlockData_T_85; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_93 = _s1_rdBlockData_T_92 | _s1_rdBlockData_T_86; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_94 = _s1_rdBlockData_T_93 | _s1_rdBlockData_T_87; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_95 = _s1_rdBlockData_T_94 | _s1_rdBlockData_T_88; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_96 = _s1_rdBlockData_T_95 | _s1_rdBlockData_T_89; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_5 = _s1_rdBlockData_T_96 | _s1_rdBlockData_T_90; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_98 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_99 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_100 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_101 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_102 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_103 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_104 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_105 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_106 = _s1_rdBlockData_T_98 | _s1_rdBlockData_T_99; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_107 = _s1_rdBlockData_T_106 | _s1_rdBlockData_T_100; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_108 = _s1_rdBlockData_T_107 | _s1_rdBlockData_T_101; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_109 = _s1_rdBlockData_T_108 | _s1_rdBlockData_T_102; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_110 = _s1_rdBlockData_T_109 | _s1_rdBlockData_T_103; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_111 = _s1_rdBlockData_T_110 | _s1_rdBlockData_T_104; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_6 = _s1_rdBlockData_T_111 | _s1_rdBlockData_T_105; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_113 = s1_info_dirInfo_chosenWay[0] ? s1_info_rdData_0_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_114 = s1_info_dirInfo_chosenWay[1] ? s1_info_rdData_1_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_115 = s1_info_dirInfo_chosenWay[2] ? s1_info_rdData_2_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_116 = s1_info_dirInfo_chosenWay[3] ? s1_info_rdData_3_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_117 = s1_info_dirInfo_chosenWay[4] ? s1_info_rdData_4_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_118 = s1_info_dirInfo_chosenWay[5] ? s1_info_rdData_5_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_119 = s1_info_dirInfo_chosenWay[6] ? s1_info_rdData_6_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_120 = s1_info_dirInfo_chosenWay[7] ? s1_info_rdData_7_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_121 = _s1_rdBlockData_T_113 | _s1_rdBlockData_T_114; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_122 = _s1_rdBlockData_T_121 | _s1_rdBlockData_T_115; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_123 = _s1_rdBlockData_T_122 | _s1_rdBlockData_T_116; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_124 = _s1_rdBlockData_T_123 | _s1_rdBlockData_T_117; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_125 = _s1_rdBlockData_T_124 | _s1_rdBlockData_T_118; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_126 = _s1_rdBlockData_T_125 | _s1_rdBlockData_T_119; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_7 = _s1_rdBlockData_T_126 | _s1_rdBlockData_T_120; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_8 = s1_blockSel[0] ? s1_rdBlockData_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_9 = s1_blockSel[1] ? s1_rdBlockData_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_10 = s1_blockSel[2] ? s1_rdBlockData_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_11 = s1_blockSel[3] ? s1_rdBlockData_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_12 = s1_blockSel[4] ? s1_rdBlockData_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_13 = s1_blockSel[5] ? s1_rdBlockData_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_14 = s1_blockSel[6] ? s1_rdBlockData_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_15 = s1_blockSel[7] ? s1_rdBlockData_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_16 = _s1_rdHitData_T_8 | _s1_rdHitData_T_9; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_17 = _s1_rdHitData_T_16 | _s1_rdHitData_T_10; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_18 = _s1_rdHitData_T_17 | _s1_rdHitData_T_11; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_19 = _s1_rdHitData_T_18 | _s1_rdHitData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_20 = _s1_rdHitData_T_19 | _s1_rdHitData_T_13; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdHitData_T_21 = _s1_rdHitData_T_20 | _s1_rdHitData_T_14; // @[Mux.scala 27:73]
  wire [31:0] s1_rdHitData = _s1_rdHitData_T_21 | _s1_rdHitData_T_15; // @[Mux.scala 27:73]
  wire  _GEN_79 = s1_full & s1_fire ? 1'h0 : s1_full; // @[ICache.scala 112:26 122:{35,45}]
  wire  _GEN_80 = s0_fire | _GEN_79; // @[ICache.scala 121:{20,30}]
  wire [1:0] _s1_bypassIdx_T = {bypassVec_1,bypassVec_0}; // @[Cat.scala 33:92]
  wire  s1_bypassIdx = _s1_bypassIdx_T[1]; // @[CircuitMath.scala 28:8]
  wire [31:0] _GEN_81 = refillBuffer_io_read_cacheLineData_0_0; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_82 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_0 : _GEN_81; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_8 = s1_blockSel[0] ? _GEN_82 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_83 = refillBuffer_io_read_cacheLineData_0_1; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_84 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_1 : _GEN_83; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_9 = s1_blockSel[1] ? _GEN_84 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_85 = refillBuffer_io_read_cacheLineData_0_2; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_86 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_2 : _GEN_85; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_10 = s1_blockSel[2] ? _GEN_86 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_87 = refillBuffer_io_read_cacheLineData_0_3; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_88 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_3 : _GEN_87; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_11 = s1_blockSel[3] ? _GEN_88 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_89 = refillBuffer_io_read_cacheLineData_0_4; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_90 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_4 : _GEN_89; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_12 = s1_blockSel[4] ? _GEN_90 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_91 = refillBuffer_io_read_cacheLineData_0_5; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_92 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_5 : _GEN_91; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_13 = s1_blockSel[5] ? _GEN_92 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_93 = refillBuffer_io_read_cacheLineData_0_6; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_94 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_6 : _GEN_93; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_14 = s1_blockSel[6] ? _GEN_94 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_95 = refillBuffer_io_read_cacheLineData_0_7; // @[Mux.scala 27:{73,73}]
  wire [31:0] _GEN_96 = s1_bypassIdx ? refillBuffer_io_read_cacheLineData_1_7 : _GEN_95; // @[Mux.scala 27:{73,73}]
  wire [31:0] _s1_bypassData_T_15 = s1_blockSel[7] ? _GEN_96 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_16 = _s1_bypassData_T_8 | _s1_bypassData_T_9; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_17 = _s1_bypassData_T_16 | _s1_bypassData_T_10; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_18 = _s1_bypassData_T_17 | _s1_bypassData_T_11; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_19 = _s1_bypassData_T_18 | _s1_bypassData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_20 = _s1_bypassData_T_19 | _s1_bypassData_T_13; // @[Mux.scala 27:73]
  wire [31:0] _s1_bypassData_T_21 = _s1_bypassData_T_20 | _s1_bypassData_T_14; // @[Mux.scala 27:73]
  reg [31:0] s2_addr; // @[Reg.scala 19:16]
  wire  _GEN_110 = s2_full & s2_fire ? 1'h0 : s2_full; // @[ICache.scala 144:26 153:{35,45}]
  wire  _GEN_111 = s1_fire | _GEN_110; // @[ICache.scala 152:{20,30}]
  wire  _refillBuffer_io_write_valid_T = io_tlbus_resp_ready & io_tlbus_resp_valid; // @[Decoupled.scala 51:35]
  wire  respHit = s1_info_dirInfo_hit & s1_full; // @[ICache.scala 166:39]
  wire  _respMiss_T_2 = refillPipe_io_resp_ready & refillPipe_io_resp_valid; // @[Decoupled.scala 51:35]
  wire  respMiss = _s2_valid_T & s2_full & _respMiss_T_2; // @[ICache.scala 167:47]
  wire  respBypass = s1_bypass & _s1_valid_T_2 & s1_full; // @[ICache.scala 168:56]
  wire [31:0] s1_bypassData = _s1_bypassData_T_21 | _s1_bypassData_T_15; // @[Mux.scala 27:73]
  wire [31:0] _io_read_resp_bits_data_T = s1_bypass ? s1_bypassData : refillPipe_io_resp_bits_data; // @[ICache.scala 172:40]
  wire [2:0] s2_off = s2_addr[4:2]; // @[ICache.scala 179:25]
  wire [3:0] rdThreshole = 4'h8 - 4'h4; // @[ICache.scala 181:41]
  wire [3:0] _GEN_112 = {{1'd0}, s1_info_req_addr[4:2]}; // @[ICache.scala 182:34]
  wire [3:0] _respHitSize_T_2 = 4'h8 - _GEN_112; // @[ICache.scala 182:68]
  wire [3:0] respHitSize = _GEN_112 >= rdThreshole ? _respHitSize_T_2 : 4'h4; // @[ICache.scala 182:26]
  wire [3:0] _GEN_114 = {{1'd0}, s2_off}; // @[ICache.scala 183:35]
  wire [3:0] _respMissSize_T_2 = 4'h8 - _GEN_114; // @[ICache.scala 183:69]
  wire [3:0] respMissSize = _GEN_114 >= rdThreshole ? _respMissSize_T_2 : 4'h4; // @[ICache.scala 183:27]
  wire [3:0] _io_read_resp_bits_size_T_1 = s1_info_dirInfo_hit | s1_bypass ? respHitSize : respMissSize; // @[ICache.scala 184:35]
  wire [255:0] _respHitInst_T = {s1_rdBlockData_7,s1_rdBlockData_6,s1_rdBlockData_5,s1_rdBlockData_4,s1_rdBlockData_3,
    s1_rdBlockData_2,s1_rdBlockData_1,s1_rdBlockData_0}; // @[ICache.scala 185:39]
  wire [7:0] _respHitInst_T_1 = {s1_info_req_addr[4:2], 5'h0}; // @[ICache.scala 185:57]
  wire [255:0] _respHitInst_T_2 = _respHitInst_T >> _respHitInst_T_1; // @[ICache.scala 185:46]
  wire [31:0] respHitInst_0 = _respHitInst_T_2[31:0]; // @[ICache.scala 185:108]
  wire [31:0] respHitInst_1 = _respHitInst_T_2[63:32]; // @[ICache.scala 185:108]
  wire [31:0] respHitInst_2 = _respHitInst_T_2[95:64]; // @[ICache.scala 185:108]
  wire [31:0] respHitInst_3 = _respHitInst_T_2[127:96]; // @[ICache.scala 185:108]
  wire [255:0] _respBypassInst_T = {_GEN_96,_GEN_94,_GEN_92,_GEN_90,_GEN_88,_GEN_86,_GEN_84,_GEN_82}; // @[ICache.scala 186:46]
  wire [255:0] _respBypassInst_T_2 = _respBypassInst_T >> _respHitInst_T_1; // @[ICache.scala 186:53]
  wire [31:0] respBypassInst_0 = _respBypassInst_T_2[31:0]; // @[ICache.scala 186:115]
  wire [31:0] respBypassInst_1 = _respBypassInst_T_2[63:32]; // @[ICache.scala 186:115]
  wire [31:0] respBypassInst_2 = _respBypassInst_T_2[95:64]; // @[ICache.scala 186:115]
  wire [31:0] respBypassInst_3 = _respBypassInst_T_2[127:96]; // @[ICache.scala 186:115]
  wire [255:0] _respRefillInst_T = {refillPipe_io_resp_bits_blockData_7,refillPipe_io_resp_bits_blockData_6,
    refillPipe_io_resp_bits_blockData_5,refillPipe_io_resp_bits_blockData_4,refillPipe_io_resp_bits_blockData_3,
    refillPipe_io_resp_bits_blockData_2,refillPipe_io_resp_bits_blockData_1,refillPipe_io_resp_bits_blockData_0}; // @[ICache.scala 187:61]
  wire [7:0] _respRefillInst_T_1 = {s2_off, 5'h0}; // @[ICache.scala 187:79]
  wire [255:0] _respRefillInst_T_2 = _respRefillInst_T >> _respRefillInst_T_1; // @[ICache.scala 187:68]
  wire [31:0] respRefillInst_0 = _respRefillInst_T_2[31:0]; // @[ICache.scala 187:130]
  wire [31:0] respRefillInst_1 = _respRefillInst_T_2[63:32]; // @[ICache.scala 187:130]
  wire [31:0] respRefillInst_2 = _respRefillInst_T_2[95:64]; // @[ICache.scala 187:130]
  wire [31:0] respRefillInst_3 = _respRefillInst_T_2[127:96]; // @[ICache.scala 187:130]
  wire [31:0] _io_read_resp_bits_inst_0_T = s1_bypass ? respBypassInst_0 : respRefillInst_0; // @[ICache.scala 191:48]
  wire [31:0] _io_read_resp_bits_inst_1_T = s1_bypass ? respBypassInst_1 : respRefillInst_1; // @[ICache.scala 191:48]
  wire [31:0] _io_read_resp_bits_inst_2_T = s1_bypass ? respBypassInst_2 : respRefillInst_2; // @[ICache.scala 191:48]
  wire [31:0] _io_read_resp_bits_inst_3_T = s1_bypass ? respBypassInst_3 : respRefillInst_3; // @[ICache.scala 191:48]
  reg [63:0] c; // @[util.scala 162:24]
  wire [63:0] _c_T_1 = c + 64'h1; // @[util.scala 163:16]
  wire [127:0] _T_7 = {io_read_resp_bits_inst_3,io_read_resp_bits_inst_2,io_read_resp_bits_inst_1,
    io_read_resp_bits_inst_0}; // @[ICache.scala 205:152]
  reg [63:0] c_1; // @[util.scala 162:24]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[util.scala 163:16]
  DataBankArray db ( // @[ICache.scala 56:20]
    .clock(db_clock),
    .reset(db_reset),
    .io_read_req_ready(db_io_read_req_ready),
    .io_read_req_valid(db_io_read_req_valid),
    .io_read_req_bits_set(db_io_read_req_bits_set),
    .io_read_resp_0_0(db_io_read_resp_0_0),
    .io_read_resp_0_1(db_io_read_resp_0_1),
    .io_read_resp_0_2(db_io_read_resp_0_2),
    .io_read_resp_0_3(db_io_read_resp_0_3),
    .io_read_resp_0_4(db_io_read_resp_0_4),
    .io_read_resp_0_5(db_io_read_resp_0_5),
    .io_read_resp_0_6(db_io_read_resp_0_6),
    .io_read_resp_0_7(db_io_read_resp_0_7),
    .io_read_resp_1_0(db_io_read_resp_1_0),
    .io_read_resp_1_1(db_io_read_resp_1_1),
    .io_read_resp_1_2(db_io_read_resp_1_2),
    .io_read_resp_1_3(db_io_read_resp_1_3),
    .io_read_resp_1_4(db_io_read_resp_1_4),
    .io_read_resp_1_5(db_io_read_resp_1_5),
    .io_read_resp_1_6(db_io_read_resp_1_6),
    .io_read_resp_1_7(db_io_read_resp_1_7),
    .io_read_resp_2_0(db_io_read_resp_2_0),
    .io_read_resp_2_1(db_io_read_resp_2_1),
    .io_read_resp_2_2(db_io_read_resp_2_2),
    .io_read_resp_2_3(db_io_read_resp_2_3),
    .io_read_resp_2_4(db_io_read_resp_2_4),
    .io_read_resp_2_5(db_io_read_resp_2_5),
    .io_read_resp_2_6(db_io_read_resp_2_6),
    .io_read_resp_2_7(db_io_read_resp_2_7),
    .io_read_resp_3_0(db_io_read_resp_3_0),
    .io_read_resp_3_1(db_io_read_resp_3_1),
    .io_read_resp_3_2(db_io_read_resp_3_2),
    .io_read_resp_3_3(db_io_read_resp_3_3),
    .io_read_resp_3_4(db_io_read_resp_3_4),
    .io_read_resp_3_5(db_io_read_resp_3_5),
    .io_read_resp_3_6(db_io_read_resp_3_6),
    .io_read_resp_3_7(db_io_read_resp_3_7),
    .io_read_resp_4_0(db_io_read_resp_4_0),
    .io_read_resp_4_1(db_io_read_resp_4_1),
    .io_read_resp_4_2(db_io_read_resp_4_2),
    .io_read_resp_4_3(db_io_read_resp_4_3),
    .io_read_resp_4_4(db_io_read_resp_4_4),
    .io_read_resp_4_5(db_io_read_resp_4_5),
    .io_read_resp_4_6(db_io_read_resp_4_6),
    .io_read_resp_4_7(db_io_read_resp_4_7),
    .io_read_resp_5_0(db_io_read_resp_5_0),
    .io_read_resp_5_1(db_io_read_resp_5_1),
    .io_read_resp_5_2(db_io_read_resp_5_2),
    .io_read_resp_5_3(db_io_read_resp_5_3),
    .io_read_resp_5_4(db_io_read_resp_5_4),
    .io_read_resp_5_5(db_io_read_resp_5_5),
    .io_read_resp_5_6(db_io_read_resp_5_6),
    .io_read_resp_5_7(db_io_read_resp_5_7),
    .io_read_resp_6_0(db_io_read_resp_6_0),
    .io_read_resp_6_1(db_io_read_resp_6_1),
    .io_read_resp_6_2(db_io_read_resp_6_2),
    .io_read_resp_6_3(db_io_read_resp_6_3),
    .io_read_resp_6_4(db_io_read_resp_6_4),
    .io_read_resp_6_5(db_io_read_resp_6_5),
    .io_read_resp_6_6(db_io_read_resp_6_6),
    .io_read_resp_6_7(db_io_read_resp_6_7),
    .io_read_resp_7_0(db_io_read_resp_7_0),
    .io_read_resp_7_1(db_io_read_resp_7_1),
    .io_read_resp_7_2(db_io_read_resp_7_2),
    .io_read_resp_7_3(db_io_read_resp_7_3),
    .io_read_resp_7_4(db_io_read_resp_7_4),
    .io_read_resp_7_5(db_io_read_resp_7_5),
    .io_read_resp_7_6(db_io_read_resp_7_6),
    .io_read_resp_7_7(db_io_read_resp_7_7),
    .io_write_req_ready(db_io_write_req_ready),
    .io_write_req_valid(db_io_write_req_valid),
    .io_write_req_bits_set(db_io_write_req_bits_set),
    .io_write_req_bits_data_0(db_io_write_req_bits_data_0),
    .io_write_req_bits_data_1(db_io_write_req_bits_data_1),
    .io_write_req_bits_data_2(db_io_write_req_bits_data_2),
    .io_write_req_bits_data_3(db_io_write_req_bits_data_3),
    .io_write_req_bits_data_4(db_io_write_req_bits_data_4),
    .io_write_req_bits_data_5(db_io_write_req_bits_data_5),
    .io_write_req_bits_data_6(db_io_write_req_bits_data_6),
    .io_write_req_bits_data_7(db_io_write_req_bits_data_7),
    .io_write_req_bits_blockMask(db_io_write_req_bits_blockMask),
    .io_write_req_bits_way(db_io_write_req_bits_way)
  );
  DCacheDirectory dir ( // @[ICache.scala 57:21]
    .clock(dir_clock),
    .reset(dir_reset),
    .io_read_req_ready(dir_io_read_req_ready),
    .io_read_req_valid(dir_io_read_req_valid),
    .io_read_req_bits_addr(dir_io_read_req_bits_addr),
    .io_read_resp_bits_hit(dir_io_read_resp_bits_hit),
    .io_read_resp_bits_chosenWay(dir_io_read_resp_bits_chosenWay),
    .io_write_req_ready(dir_io_write_req_ready),
    .io_write_req_valid(dir_io_write_req_valid),
    .io_write_req_bits_addr(dir_io_write_req_bits_addr),
    .io_write_req_bits_way(dir_io_write_req_bits_way)
  );
  RefillPipe refillPipe ( // @[ICache.scala 58:28]
    .clock(refillPipe_clock),
    .reset(refillPipe_reset),
    .io_req_ready(refillPipe_io_req_ready),
    .io_req_valid(refillPipe_io_req_valid),
    .io_req_bits_addr(refillPipe_io_req_bits_addr),
    .io_req_bits_chosenWay(refillPipe_io_req_bits_chosenWay),
    .io_resp_ready(refillPipe_io_resp_ready),
    .io_resp_valid(refillPipe_io_resp_valid),
    .io_resp_bits_data(refillPipe_io_resp_bits_data),
    .io_resp_bits_blockData_0(refillPipe_io_resp_bits_blockData_0),
    .io_resp_bits_blockData_1(refillPipe_io_resp_bits_blockData_1),
    .io_resp_bits_blockData_2(refillPipe_io_resp_bits_blockData_2),
    .io_resp_bits_blockData_3(refillPipe_io_resp_bits_blockData_3),
    .io_resp_bits_blockData_4(refillPipe_io_resp_bits_blockData_4),
    .io_resp_bits_blockData_5(refillPipe_io_resp_bits_blockData_5),
    .io_resp_bits_blockData_6(refillPipe_io_resp_bits_blockData_6),
    .io_resp_bits_blockData_7(refillPipe_io_resp_bits_blockData_7),
    .io_tlbus_req_ready(refillPipe_io_tlbus_req_ready),
    .io_tlbus_req_valid(refillPipe_io_tlbus_req_valid),
    .io_tlbus_req_bits_size(refillPipe_io_tlbus_req_bits_size),
    .io_tlbus_req_bits_address(refillPipe_io_tlbus_req_bits_address),
    .io_tlbus_resp_ready(refillPipe_io_tlbus_resp_ready),
    .io_tlbus_resp_valid(refillPipe_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(refillPipe_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(refillPipe_io_tlbus_resp_bits_data),
    .io_dirWrite_req_valid(refillPipe_io_dirWrite_req_valid),
    .io_dirWrite_req_bits_addr(refillPipe_io_dirWrite_req_bits_addr),
    .io_dirWrite_req_bits_way(refillPipe_io_dirWrite_req_bits_way),
    .io_dataWrite_req_valid(refillPipe_io_dataWrite_req_valid),
    .io_dataWrite_req_bits_set(refillPipe_io_dataWrite_req_bits_set),
    .io_dataWrite_req_bits_data_0(refillPipe_io_dataWrite_req_bits_data_0),
    .io_dataWrite_req_bits_data_1(refillPipe_io_dataWrite_req_bits_data_1),
    .io_dataWrite_req_bits_data_2(refillPipe_io_dataWrite_req_bits_data_2),
    .io_dataWrite_req_bits_data_3(refillPipe_io_dataWrite_req_bits_data_3),
    .io_dataWrite_req_bits_data_4(refillPipe_io_dataWrite_req_bits_data_4),
    .io_dataWrite_req_bits_data_5(refillPipe_io_dataWrite_req_bits_data_5),
    .io_dataWrite_req_bits_data_6(refillPipe_io_dataWrite_req_bits_data_6),
    .io_dataWrite_req_bits_data_7(refillPipe_io_dataWrite_req_bits_data_7),
    .io_dataWrite_req_bits_blockMask(refillPipe_io_dataWrite_req_bits_blockMask),
    .io_dataWrite_req_bits_way(refillPipe_io_dataWrite_req_bits_way)
  );
  RefillBuffer refillBuffer ( // @[ICache.scala 65:30]
    .clock(refillBuffer_clock),
    .reset(refillBuffer_reset),
    .io_write_valid(refillBuffer_io_write_valid),
    .io_write_bits_cacheLineAddr(refillBuffer_io_write_bits_cacheLineAddr),
    .io_write_bits_data(refillBuffer_io_write_bits_data),
    .io_read_cacheLineAddr_0(refillBuffer_io_read_cacheLineAddr_0),
    .io_read_cacheLineAddr_1(refillBuffer_io_read_cacheLineAddr_1),
    .io_read_cacheLineData_0_0(refillBuffer_io_read_cacheLineData_0_0),
    .io_read_cacheLineData_0_1(refillBuffer_io_read_cacheLineData_0_1),
    .io_read_cacheLineData_0_2(refillBuffer_io_read_cacheLineData_0_2),
    .io_read_cacheLineData_0_3(refillBuffer_io_read_cacheLineData_0_3),
    .io_read_cacheLineData_0_4(refillBuffer_io_read_cacheLineData_0_4),
    .io_read_cacheLineData_0_5(refillBuffer_io_read_cacheLineData_0_5),
    .io_read_cacheLineData_0_6(refillBuffer_io_read_cacheLineData_0_6),
    .io_read_cacheLineData_0_7(refillBuffer_io_read_cacheLineData_0_7),
    .io_read_cacheLineData_1_0(refillBuffer_io_read_cacheLineData_1_0),
    .io_read_cacheLineData_1_1(refillBuffer_io_read_cacheLineData_1_1),
    .io_read_cacheLineData_1_2(refillBuffer_io_read_cacheLineData_1_2),
    .io_read_cacheLineData_1_3(refillBuffer_io_read_cacheLineData_1_3),
    .io_read_cacheLineData_1_4(refillBuffer_io_read_cacheLineData_1_4),
    .io_read_cacheLineData_1_5(refillBuffer_io_read_cacheLineData_1_5),
    .io_read_cacheLineData_1_6(refillBuffer_io_read_cacheLineData_1_6),
    .io_read_cacheLineData_1_7(refillBuffer_io_read_cacheLineData_1_7),
    .io_read_valids_0(refillBuffer_io_read_valids_0),
    .io_read_valids_1(refillBuffer_io_read_valids_1)
  );
  assign io_read_req_ready = ~s0_full | s0_fire; // @[ICache.scala 80:35]
  assign io_read_resp_valid = respHit | respMiss | respBypass; // @[ICache.scala 169:48]
  assign io_read_resp_bits_data = s1_info_dirInfo_hit ? s1_rdHitData : _io_read_resp_bits_data_T; // @[ICache.scala 170:34]
  assign io_read_resp_bits_inst_0 = s1_info_dirInfo_hit ? respHitInst_0 : _io_read_resp_bits_inst_0_T; // @[ICache.scala 189:41]
  assign io_read_resp_bits_inst_1 = s1_info_dirInfo_hit ? respHitInst_1 : _io_read_resp_bits_inst_1_T; // @[ICache.scala 189:41]
  assign io_read_resp_bits_inst_2 = s1_info_dirInfo_hit ? respHitInst_2 : _io_read_resp_bits_inst_2_T; // @[ICache.scala 189:41]
  assign io_read_resp_bits_inst_3 = s1_info_dirInfo_hit ? respHitInst_3 : _io_read_resp_bits_inst_3_T; // @[ICache.scala 189:41]
  assign io_read_resp_bits_size = _io_read_resp_bits_size_T_1[2:0]; // @[ICache.scala 184:28]
  assign io_tlbus_req_valid = refillPipe_io_tlbus_req_valid; // @[ICache.scala 63:25]
  assign io_tlbus_req_bits_address = refillPipe_io_tlbus_req_bits_address; // @[ICache.scala 63:25]
  assign io_tlbus_resp_ready = 1'h1; // @[ICache.scala 201:25]
  assign db_clock = clock;
  assign db_reset = reset;
  assign db_io_read_req_valid = s0_latch | s0_full; // @[ICache.scala 85:38]
  assign db_io_read_req_bits_set = _GEN_0[11:5]; // @[Parameters.scala 50:11]
  assign db_io_write_req_valid = refillPipe_io_dataWrite_req_valid; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_set = refillPipe_io_dataWrite_req_bits_set; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_data_0 = refillPipe_io_dataWrite_req_bits_data_0; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_data_1 = refillPipe_io_dataWrite_req_bits_data_1; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_data_2 = refillPipe_io_dataWrite_req_bits_data_2; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_data_3 = refillPipe_io_dataWrite_req_bits_data_3; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_data_4 = refillPipe_io_dataWrite_req_bits_data_4; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_data_5 = refillPipe_io_dataWrite_req_bits_data_5; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_data_6 = refillPipe_io_dataWrite_req_bits_data_6; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_data_7 = refillPipe_io_dataWrite_req_bits_data_7; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_blockMask = refillPipe_io_dataWrite_req_bits_blockMask; // @[ICache.scala 61:33]
  assign db_io_write_req_bits_way = refillPipe_io_dataWrite_req_bits_way; // @[ICache.scala 61:33]
  assign dir_clock = clock;
  assign dir_reset = reset;
  assign dir_io_read_req_valid = s0_latch | s0_full; // @[ICache.scala 88:39]
  assign dir_io_read_req_bits_addr = s0_latch ? io_read_req_bits_addr : s0_req_r_addr; // @[ICache.scala 78:21]
  assign dir_io_write_req_valid = refillPipe_io_dirWrite_req_valid; // @[ICache.scala 62:32]
  assign dir_io_write_req_bits_addr = refillPipe_io_dirWrite_req_bits_addr; // @[ICache.scala 62:32]
  assign dir_io_write_req_bits_way = refillPipe_io_dirWrite_req_bits_way; // @[ICache.scala 62:32]
  assign refillPipe_clock = clock;
  assign refillPipe_reset = reset;
  assign refillPipe_io_req_valid = _s1_valid_T_2 & s1_full & _s1_valid_T_5; // @[ICache.scala 132:64]
  assign refillPipe_io_req_bits_addr = s1_info_req_addr; // @[ICache.scala 133:33]
  assign refillPipe_io_req_bits_chosenWay = s1_info_dirInfo_chosenWay; // @[ICache.scala 134:38]
  assign refillPipe_io_resp_ready = 1'h1; // @[ICache.scala 199:30]
  assign refillPipe_io_tlbus_req_ready = io_tlbus_req_ready; // @[ICache.scala 63:25]
  assign refillPipe_io_tlbus_resp_valid = io_tlbus_resp_valid; // @[ICache.scala 63:25]
  assign refillPipe_io_tlbus_resp_bits_opcode = io_tlbus_resp_bits_opcode; // @[ICache.scala 63:25]
  assign refillPipe_io_tlbus_resp_bits_data = io_tlbus_resp_bits_data; // @[ICache.scala 63:25]
  assign refillBuffer_clock = clock;
  assign refillBuffer_reset = reset;
  assign refillBuffer_io_write_valid = _refillBuffer_io_write_valid_T & io_tlbus_resp_bits_opcode == 3'h1; // @[ICache.scala 156:55]
  assign refillBuffer_io_write_bits_cacheLineAddr = s2_addr; // @[ICache.scala 158:46]
  assign refillBuffer_io_write_bits_data = io_tlbus_resp_bits_data; // @[ICache.scala 157:37]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 75:26]
      s0_full <= 1'h0; // @[ICache.scala 75:26]
    end else begin
      s0_full <= _GEN_2;
    end
    if (reset) begin // @[ICache.scala 112:26]
      s1_full <= 1'h0; // @[ICache.scala 112:26]
    end else begin
      s1_full <= _GEN_80;
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_dirInfo_hit <= s0_info_dirInfo_hit; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      if (s0_latch) begin // @[Reg.scala 20:18]
        s1_info_req_addr <= io_read_req_bits_addr; // @[Reg.scala 20:22]
      end else begin
        s1_info_req_addr <= s0_req_r_addr; // @[Reg.scala 19:16]
      end
    end
    if (reset) begin // @[ICache.scala 144:26]
      s2_full <= 1'h0; // @[ICache.scala 144:26]
    end else begin
      s2_full <= _GEN_111;
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_dirInfo_hit <= s1_info_dirInfo_hit; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_bypass <= s1_bypass; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_req_r_addr <= io_read_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_dirInfo_chosenWay <= s0_info_dirInfo_chosenWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_0 <= s0_info_rdData_0_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_1 <= s0_info_rdData_0_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_2 <= s0_info_rdData_0_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_3 <= s0_info_rdData_0_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_4 <= s0_info_rdData_0_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_5 <= s0_info_rdData_0_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_6 <= s0_info_rdData_0_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_0_7 <= s0_info_rdData_0_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_0 <= s0_info_rdData_1_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_1 <= s0_info_rdData_1_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_2 <= s0_info_rdData_1_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_3 <= s0_info_rdData_1_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_4 <= s0_info_rdData_1_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_5 <= s0_info_rdData_1_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_6 <= s0_info_rdData_1_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_1_7 <= s0_info_rdData_1_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_0 <= s0_info_rdData_2_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_1 <= s0_info_rdData_2_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_2 <= s0_info_rdData_2_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_3 <= s0_info_rdData_2_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_4 <= s0_info_rdData_2_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_5 <= s0_info_rdData_2_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_6 <= s0_info_rdData_2_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_2_7 <= s0_info_rdData_2_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_0 <= s0_info_rdData_3_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_1 <= s0_info_rdData_3_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_2 <= s0_info_rdData_3_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_3 <= s0_info_rdData_3_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_4 <= s0_info_rdData_3_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_5 <= s0_info_rdData_3_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_6 <= s0_info_rdData_3_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_3_7 <= s0_info_rdData_3_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_0 <= s0_info_rdData_4_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_1 <= s0_info_rdData_4_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_2 <= s0_info_rdData_4_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_3 <= s0_info_rdData_4_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_4 <= s0_info_rdData_4_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_5 <= s0_info_rdData_4_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_6 <= s0_info_rdData_4_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_4_7 <= s0_info_rdData_4_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_0 <= s0_info_rdData_5_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_1 <= s0_info_rdData_5_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_2 <= s0_info_rdData_5_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_3 <= s0_info_rdData_5_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_4 <= s0_info_rdData_5_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_5 <= s0_info_rdData_5_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_6 <= s0_info_rdData_5_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_5_7 <= s0_info_rdData_5_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_0 <= s0_info_rdData_6_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_1 <= s0_info_rdData_6_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_2 <= s0_info_rdData_6_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_3 <= s0_info_rdData_6_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_4 <= s0_info_rdData_6_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_5 <= s0_info_rdData_6_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_6 <= s0_info_rdData_6_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_6_7 <= s0_info_rdData_6_7; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_0 <= s0_info_rdData_7_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_1 <= s0_info_rdData_7_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_2 <= s0_info_rdData_7_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_3 <= s0_info_rdData_7_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_4 <= s0_info_rdData_7_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_5 <= s0_info_rdData_7_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_6 <= s0_info_rdData_7_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_info_rdData_7_7 <= s0_info_rdData_7_7; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_addr <= s1_info_req_addr; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[util.scala 162:24]
      c <= 64'h0; // @[util.scala 162:24]
    end else begin
      c <= _c_T_1; // @[util.scala 163:11]
    end
    if (reset) begin // @[util.scala 162:24]
      c_1 <= 64'h0; // @[util.scala 162:24]
    end else begin
      c_1 <= _c_T_3; // @[util.scala 163:11]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s0_latch & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [ICache] read req ==> addr: 0x%x\n",c,io_read_req_bits_addr); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_read_resp_valid & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [ICache] read resp <== data: 0x%x  inst:0x%x\n",c_1,
            io_read_resp_bits_data,_T_7); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s1_full = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s1_info_dirInfo_hit = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s1_info_req_addr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  s2_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s2_dirInfo_hit = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s2_bypass = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s0_req_r_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  s1_info_dirInfo_chosenWay = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  s1_info_rdData_0_0 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  s1_info_rdData_0_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  s1_info_rdData_0_2 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  s1_info_rdData_0_3 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  s1_info_rdData_0_4 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  s1_info_rdData_0_5 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  s1_info_rdData_0_6 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  s1_info_rdData_0_7 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  s1_info_rdData_1_0 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  s1_info_rdData_1_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  s1_info_rdData_1_2 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  s1_info_rdData_1_3 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  s1_info_rdData_1_4 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  s1_info_rdData_1_5 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  s1_info_rdData_1_6 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  s1_info_rdData_1_7 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  s1_info_rdData_2_0 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  s1_info_rdData_2_1 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  s1_info_rdData_2_2 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  s1_info_rdData_2_3 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  s1_info_rdData_2_4 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  s1_info_rdData_2_5 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  s1_info_rdData_2_6 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  s1_info_rdData_2_7 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  s1_info_rdData_3_0 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  s1_info_rdData_3_1 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  s1_info_rdData_3_2 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  s1_info_rdData_3_3 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  s1_info_rdData_3_4 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  s1_info_rdData_3_5 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  s1_info_rdData_3_6 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  s1_info_rdData_3_7 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  s1_info_rdData_4_0 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  s1_info_rdData_4_1 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  s1_info_rdData_4_2 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  s1_info_rdData_4_3 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  s1_info_rdData_4_4 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  s1_info_rdData_4_5 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  s1_info_rdData_4_6 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  s1_info_rdData_4_7 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  s1_info_rdData_5_0 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  s1_info_rdData_5_1 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  s1_info_rdData_5_2 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  s1_info_rdData_5_3 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  s1_info_rdData_5_4 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  s1_info_rdData_5_5 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  s1_info_rdData_5_6 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  s1_info_rdData_5_7 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  s1_info_rdData_6_0 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  s1_info_rdData_6_1 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  s1_info_rdData_6_2 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  s1_info_rdData_6_3 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  s1_info_rdData_6_4 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  s1_info_rdData_6_5 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  s1_info_rdData_6_6 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  s1_info_rdData_6_7 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  s1_info_rdData_7_0 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  s1_info_rdData_7_1 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  s1_info_rdData_7_2 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  s1_info_rdData_7_3 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  s1_info_rdData_7_4 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  s1_info_rdData_7_5 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  s1_info_rdData_7_6 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  s1_info_rdData_7_7 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  s2_addr = _RAND_73[31:0];
  _RAND_74 = {2{`RANDOM}};
  c = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  c_1 = _RAND_75[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Fetch_1(
  input          clock,
  input          reset,
  input          io_in_start,
  input          io_in_execute_bits_brTaken,
  input  [31:0]  io_in_execute_bits_targetAddr,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_pcNext4,
  output         io_out_bits_instState_commit,
  output [31:0]  io_out_bits_instState_pc,
  output [31:0]  io_out_bits_instState_inst,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [31:0]  io_tlbus_req_bits_address,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data,
  input  [31:0]  io_trapVec,
  input  [31:0]  io_mepc,
  input          io_excp_valid,
  input          io_excp_bits_isMret
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  icache_clock; // @[1_Fetch.scala 151:24]
  wire  icache_reset; // @[1_Fetch.scala 151:24]
  wire  icache_io_read_req_ready; // @[1_Fetch.scala 151:24]
  wire  icache_io_read_req_valid; // @[1_Fetch.scala 151:24]
  wire [31:0] icache_io_read_req_bits_addr; // @[1_Fetch.scala 151:24]
  wire  icache_io_read_resp_ready; // @[1_Fetch.scala 151:24]
  wire  icache_io_read_resp_valid; // @[1_Fetch.scala 151:24]
  wire [31:0] icache_io_read_resp_bits_data; // @[1_Fetch.scala 151:24]
  wire [31:0] icache_io_read_resp_bits_inst_0; // @[1_Fetch.scala 151:24]
  wire [31:0] icache_io_read_resp_bits_inst_1; // @[1_Fetch.scala 151:24]
  wire [31:0] icache_io_read_resp_bits_inst_2; // @[1_Fetch.scala 151:24]
  wire [31:0] icache_io_read_resp_bits_inst_3; // @[1_Fetch.scala 151:24]
  wire [2:0] icache_io_read_resp_bits_size; // @[1_Fetch.scala 151:24]
  wire  icache_io_tlbus_req_ready; // @[1_Fetch.scala 151:24]
  wire  icache_io_tlbus_req_valid; // @[1_Fetch.scala 151:24]
  wire [31:0] icache_io_tlbus_req_bits_address; // @[1_Fetch.scala 151:24]
  wire  icache_io_tlbus_resp_ready; // @[1_Fetch.scala 151:24]
  wire  icache_io_tlbus_resp_valid; // @[1_Fetch.scala 151:24]
  wire [2:0] icache_io_tlbus_resp_bits_opcode; // @[1_Fetch.scala 151:24]
  wire [127:0] icache_io_tlbus_resp_bits_data; // @[1_Fetch.scala 151:24]
  reg [31:0] pcReg; // @[1_Fetch.scala 137:34]
  wire [31:0] pcNext4 = pcReg + 32'h4; // @[1_Fetch.scala 139:33]
  wire [31:0] _branchAddr_1_T = io_excp_bits_isMret ? io_mepc : io_trapVec; // @[1_Fetch.scala 142:24]
  wire [31:0] _branchAddr_1_T_1 = io_in_execute_bits_brTaken ? io_in_execute_bits_targetAddr : pcReg; // @[1_Fetch.scala 146:24]
  wire [31:0] branchAddr_1 = io_excp_valid ? _branchAddr_1_T : _branchAddr_1_T_1; // @[1_Fetch.scala 141:27]
  wire  hasBranch_1 = io_excp_valid | io_in_execute_bits_brTaken; // @[1_Fetch.scala 164:37]
  wire  _hasBranch_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire  _hasBranch_T_1 = ~io_in_start; // @[1_Fetch.scala 165:62]
  wire  _hasBranch_T_2 = _hasBranch_T | ~io_in_start; // @[1_Fetch.scala 165:59]
  reg  hasBranch_holdReg; // @[Reg.scala 19:16]
  wire  _GEN_0 = hasBranch_1 | hasBranch_holdReg; // @[Reg.scala 19:16 20:{18,22}]
  wire  hasBranch = hasBranch_1 | hasBranch_holdReg; // @[util.scala 26:12]
  reg [31:0] branchAddr_holdReg; // @[Reg.scala 19:16]
  wire [31:0] _GEN_2 = hasBranch_1 ? branchAddr_1 : branchAddr_holdReg; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] pcNext = _GEN_0 ? _GEN_2 : pcNext4; // @[1_Fetch.scala 169:18]
  wire  commit = io_out_ready & ~_GEN_0; // @[1_Fetch.scala 177:50]
  wire  _lastInstValid_T = icache_io_read_resp_ready & icache_io_read_resp_valid; // @[Decoupled.scala 51:35]
  reg  lastInstValid_holdReg; // @[Reg.scala 19:16]
  wire  _GEN_4 = _lastInstValid_T | lastInstValid_holdReg; // @[Reg.scala 19:16 20:{18,22}]
  wire  lastInstValid = _lastInstValid_T | lastInstValid_holdReg; // @[util.scala 26:12]
  wire  _firstFire_T = icache_io_read_req_ready & icache_io_read_req_valid; // @[Decoupled.scala 51:35]
  reg  firstFire; // @[Reg.scala 35:20]
  wire  _GEN_6 = _firstFire_T ? 1'h0 : firstFire; // @[Reg.scala 36:18 35:20 36:22]
  wire  preFetchInst = firstFire & pcReg == 32'h0 | ~firstFire & _hasBranch_T; // @[1_Fetch.scala 183:59]
  reg [31:0] inst_r; // @[Reg.scala 19:16]
  wire [31:0] _GEN_7 = _lastInstValid_T ? icache_io_read_resp_bits_data : inst_r; // @[Reg.scala 19:16 20:{18,22}]
  ICache icache ( // @[1_Fetch.scala 151:24]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_read_req_ready(icache_io_read_req_ready),
    .io_read_req_valid(icache_io_read_req_valid),
    .io_read_req_bits_addr(icache_io_read_req_bits_addr),
    .io_read_resp_ready(icache_io_read_resp_ready),
    .io_read_resp_valid(icache_io_read_resp_valid),
    .io_read_resp_bits_data(icache_io_read_resp_bits_data),
    .io_read_resp_bits_inst_0(icache_io_read_resp_bits_inst_0),
    .io_read_resp_bits_inst_1(icache_io_read_resp_bits_inst_1),
    .io_read_resp_bits_inst_2(icache_io_read_resp_bits_inst_2),
    .io_read_resp_bits_inst_3(icache_io_read_resp_bits_inst_3),
    .io_read_resp_bits_size(icache_io_read_resp_bits_size),
    .io_tlbus_req_ready(icache_io_tlbus_req_ready),
    .io_tlbus_req_valid(icache_io_tlbus_req_valid),
    .io_tlbus_req_bits_address(icache_io_tlbus_req_bits_address),
    .io_tlbus_resp_ready(icache_io_tlbus_resp_ready),
    .io_tlbus_resp_valid(icache_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(icache_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(icache_io_tlbus_resp_bits_data)
  );
  assign io_out_valid = io_in_start & icache_io_read_req_ready & _GEN_4; // @[1_Fetch.scala 206:71]
  assign io_out_bits_pcNext4 = pcReg + 32'h4; // @[1_Fetch.scala 139:33]
  assign io_out_bits_instState_commit = io_out_ready & ~_GEN_0; // @[1_Fetch.scala 177:50]
  assign io_out_bits_instState_pc = pcReg; // @[1_Fetch.scala 201:19 198:34]
  assign io_out_bits_instState_inst = commit ? _GEN_7 : 32'h13; // @[1_Fetch.scala 199:40]
  assign io_tlbus_req_valid = icache_io_tlbus_req_valid; // @[1_Fetch.scala 185:21]
  assign io_tlbus_req_bits_address = icache_io_tlbus_req_bits_address; // @[1_Fetch.scala 185:21]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_read_req_valid = io_in_start & preFetchInst; // @[1_Fetch.scala 186:55]
  assign icache_io_read_req_bits_addr = _hasBranch_T ? pcNext : pcReg; // @[1_Fetch.scala 187:40]
  assign icache_io_read_resp_ready = 1'h1; // @[1_Fetch.scala 188:31]
  assign icache_io_tlbus_req_ready = io_tlbus_req_ready; // @[1_Fetch.scala 185:21]
  assign icache_io_tlbus_resp_valid = io_tlbus_resp_valid; // @[1_Fetch.scala 185:21]
  assign icache_io_tlbus_resp_bits_opcode = io_tlbus_resp_bits_opcode; // @[1_Fetch.scala 185:21]
  assign icache_io_tlbus_resp_bits_data = io_tlbus_resp_bits_data; // @[1_Fetch.scala 185:21]
  always @(posedge clock) begin
    if (reset) begin // @[1_Fetch.scala 137:34]
      pcReg <= 32'h0; // @[1_Fetch.scala 137:34]
    end else if (_hasBranch_T) begin // @[1_Fetch.scala 187:40]
      if (_GEN_0) begin // @[1_Fetch.scala 169:18]
        if (hasBranch_1) begin // @[Reg.scala 20:18]
          pcReg <= branchAddr_1; // @[Reg.scala 20:22]
        end else begin
          pcReg <= branchAddr_holdReg; // @[Reg.scala 19:16]
        end
      end else begin
        pcReg <= pcNext4;
      end
    end
    if (_hasBranch_T_2) begin // @[util.scala 25:21]
      hasBranch_holdReg <= 1'h0; // @[util.scala 25:31]
    end else begin
      hasBranch_holdReg <= _GEN_0;
    end
    if (_hasBranch_T_1) begin // @[util.scala 25:21]
      branchAddr_holdReg <= 32'h0; // @[util.scala 25:31]
    end else if (hasBranch_1) begin // @[Reg.scala 20:18]
      if (io_excp_valid) begin // @[1_Fetch.scala 141:27]
        if (io_excp_bits_isMret) begin // @[1_Fetch.scala 142:24]
          branchAddr_holdReg <= io_mepc;
        end else begin
          branchAddr_holdReg <= io_trapVec;
        end
      end else if (io_in_execute_bits_brTaken) begin // @[1_Fetch.scala 146:24]
        branchAddr_holdReg <= io_in_execute_bits_targetAddr;
      end else begin
        branchAddr_holdReg <= pcReg;
      end
    end
    if (_hasBranch_T) begin // @[util.scala 25:21]
      lastInstValid_holdReg <= 1'h0; // @[util.scala 25:31]
    end else begin
      lastInstValid_holdReg <= _GEN_4;
    end
    firstFire <= reset | _GEN_6; // @[Reg.scala 35:{20,20}]
    if (_lastInstValid_T) begin // @[Reg.scala 20:18]
      inst_r <= icache_io_read_resp_bits_data; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  hasBranch_holdReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  branchAddr_holdReg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  lastInstValid_holdReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  firstFire = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  inst_r = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decoder(
  input  [31:0] io_inst,
  output        io_out_isBranch,
  output [1:0]  io_out_resultSrc,
  output [3:0]  io_out_aluOpSel,
  output [4:0]  io_out_lsuOp,
  output [3:0]  io_out_aluSrc1,
  output [3:0]  io_out_aluSrc2,
  output [2:0]  io_out_immSrc,
  output        io_out_immSign,
  output        io_out_regWrEn,
  output [2:0]  io_out_csrOp,
  output [3:0]  io_out_excType
);
  wire [31:0] _decodeSigs_T = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_1 = 32'h3 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_3 = 32'h1003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_5 = 32'h2003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_7 = 32'h4003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_9 = 32'h5003 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_11 = 32'h13 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [31:0] _decodeSigs_T_12 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_13 = 32'h1013 == _decodeSigs_T_12; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_15 = 32'h2013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_17 = 32'h3013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_19 = 32'h4013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_21 = 32'h5013 == _decodeSigs_T_12; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_23 = 32'h40005013 == _decodeSigs_T_12; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_25 = 32'h6013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_27 = 32'h7013 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [31:0] _decodeSigs_T_28 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_29 = 32'h17 == _decodeSigs_T_28; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_31 = 32'h23 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_33 = 32'h1023 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_35 = 32'h2023 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire [31:0] _decodeSigs_T_36 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_37 = 32'h33 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_39 = 32'h40000033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_41 = 32'h1033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_43 = 32'h2033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_45 = 32'h3033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_47 = 32'h4033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_49 = 32'h5033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_51 = 32'h40005033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_53 = 32'h6033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_55 = 32'h7033 == _decodeSigs_T_36; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_57 = 32'h37 == _decodeSigs_T_28; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_59 = 32'h63 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_61 = 32'h1063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_63 = 32'h4063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_65 = 32'h5063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_67 = 32'h6063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_69 = 32'h7063 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_71 = 32'h67 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_73 = 32'h6f == _decodeSigs_T_28; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_75 = 32'hf == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_77 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_79 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_81 = 32'h30200073 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_83 = 32'h10200073 == io_inst; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_85 = 32'h1073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_87 = 32'h2073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_89 = 32'h3073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_91 = 32'h5073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_93 = 32'h6073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_95 = 32'h7073 == _decodeSigs_T; // @[Lookup.scala 31:38]
  wire  _decodeSigs_T_115 = _decodeSigs_T_57 ? 1'h0 : _decodeSigs_T_59 | (_decodeSigs_T_61 | (_decodeSigs_T_63 | (
    _decodeSigs_T_65 | (_decodeSigs_T_67 | _decodeSigs_T_69)))); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_116 = _decodeSigs_T_55 ? 1'h0 : _decodeSigs_T_115; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_117 = _decodeSigs_T_53 ? 1'h0 : _decodeSigs_T_116; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_118 = _decodeSigs_T_51 ? 1'h0 : _decodeSigs_T_117; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_119 = _decodeSigs_T_49 ? 1'h0 : _decodeSigs_T_118; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_120 = _decodeSigs_T_47 ? 1'h0 : _decodeSigs_T_119; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_121 = _decodeSigs_T_45 ? 1'h0 : _decodeSigs_T_120; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_122 = _decodeSigs_T_43 ? 1'h0 : _decodeSigs_T_121; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_123 = _decodeSigs_T_41 ? 1'h0 : _decodeSigs_T_122; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_124 = _decodeSigs_T_39 ? 1'h0 : _decodeSigs_T_123; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_125 = _decodeSigs_T_37 ? 1'h0 : _decodeSigs_T_124; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_126 = _decodeSigs_T_35 ? 1'h0 : _decodeSigs_T_125; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_127 = _decodeSigs_T_33 ? 1'h0 : _decodeSigs_T_126; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_128 = _decodeSigs_T_31 ? 1'h0 : _decodeSigs_T_127; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_129 = _decodeSigs_T_29 ? 1'h0 : _decodeSigs_T_128; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_130 = _decodeSigs_T_27 ? 1'h0 : _decodeSigs_T_129; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_131 = _decodeSigs_T_25 ? 1'h0 : _decodeSigs_T_130; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_132 = _decodeSigs_T_23 ? 1'h0 : _decodeSigs_T_131; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_133 = _decodeSigs_T_21 ? 1'h0 : _decodeSigs_T_132; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_134 = _decodeSigs_T_19 ? 1'h0 : _decodeSigs_T_133; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_135 = _decodeSigs_T_17 ? 1'h0 : _decodeSigs_T_134; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_136 = _decodeSigs_T_15 ? 1'h0 : _decodeSigs_T_135; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_137 = _decodeSigs_T_13 ? 1'h0 : _decodeSigs_T_136; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_138 = _decodeSigs_T_11 ? 1'h0 : _decodeSigs_T_137; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_139 = _decodeSigs_T_9 ? 1'h0 : _decodeSigs_T_138; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_140 = _decodeSigs_T_7 ? 1'h0 : _decodeSigs_T_139; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_141 = _decodeSigs_T_5 ? 1'h0 : _decodeSigs_T_140; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_142 = _decodeSigs_T_3 ? 1'h0 : _decodeSigs_T_141; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_143 = _decodeSigs_T_95 ? 2'h3 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_144 = _decodeSigs_T_93 ? 2'h3 : _decodeSigs_T_143; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_145 = _decodeSigs_T_91 ? 2'h3 : _decodeSigs_T_144; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_146 = _decodeSigs_T_89 ? 2'h3 : _decodeSigs_T_145; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_147 = _decodeSigs_T_87 ? 2'h3 : _decodeSigs_T_146; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_148 = _decodeSigs_T_85 ? 2'h3 : _decodeSigs_T_147; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_149 = _decodeSigs_T_83 ? 2'h0 : _decodeSigs_T_148; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_150 = _decodeSigs_T_81 ? 2'h0 : _decodeSigs_T_149; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_151 = _decodeSigs_T_79 ? 2'h0 : _decodeSigs_T_150; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_152 = _decodeSigs_T_77 ? 2'h0 : _decodeSigs_T_151; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_153 = _decodeSigs_T_75 ? 2'h0 : _decodeSigs_T_152; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_154 = _decodeSigs_T_73 ? 2'h2 : _decodeSigs_T_153; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_155 = _decodeSigs_T_71 ? 2'h2 : _decodeSigs_T_154; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_156 = _decodeSigs_T_69 ? 2'h0 : _decodeSigs_T_155; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_157 = _decodeSigs_T_67 ? 2'h0 : _decodeSigs_T_156; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_158 = _decodeSigs_T_65 ? 2'h0 : _decodeSigs_T_157; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_159 = _decodeSigs_T_63 ? 2'h0 : _decodeSigs_T_158; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_160 = _decodeSigs_T_61 ? 2'h0 : _decodeSigs_T_159; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_161 = _decodeSigs_T_59 ? 2'h0 : _decodeSigs_T_160; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_162 = _decodeSigs_T_57 ? 2'h0 : _decodeSigs_T_161; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_163 = _decodeSigs_T_55 ? 2'h0 : _decodeSigs_T_162; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_164 = _decodeSigs_T_53 ? 2'h0 : _decodeSigs_T_163; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_165 = _decodeSigs_T_51 ? 2'h0 : _decodeSigs_T_164; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_166 = _decodeSigs_T_49 ? 2'h0 : _decodeSigs_T_165; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_167 = _decodeSigs_T_47 ? 2'h0 : _decodeSigs_T_166; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_168 = _decodeSigs_T_45 ? 2'h0 : _decodeSigs_T_167; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_169 = _decodeSigs_T_43 ? 2'h0 : _decodeSigs_T_168; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_170 = _decodeSigs_T_41 ? 2'h0 : _decodeSigs_T_169; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_171 = _decodeSigs_T_39 ? 2'h0 : _decodeSigs_T_170; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_172 = _decodeSigs_T_37 ? 2'h0 : _decodeSigs_T_171; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_173 = _decodeSigs_T_35 ? 2'h0 : _decodeSigs_T_172; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_174 = _decodeSigs_T_33 ? 2'h0 : _decodeSigs_T_173; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_175 = _decodeSigs_T_31 ? 2'h0 : _decodeSigs_T_174; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_176 = _decodeSigs_T_29 ? 2'h0 : _decodeSigs_T_175; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_177 = _decodeSigs_T_27 ? 2'h0 : _decodeSigs_T_176; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_178 = _decodeSigs_T_25 ? 2'h0 : _decodeSigs_T_177; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_179 = _decodeSigs_T_23 ? 2'h0 : _decodeSigs_T_178; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_180 = _decodeSigs_T_21 ? 2'h0 : _decodeSigs_T_179; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_181 = _decodeSigs_T_19 ? 2'h0 : _decodeSigs_T_180; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_182 = _decodeSigs_T_17 ? 2'h0 : _decodeSigs_T_181; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_183 = _decodeSigs_T_15 ? 2'h0 : _decodeSigs_T_182; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_184 = _decodeSigs_T_13 ? 2'h0 : _decodeSigs_T_183; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_185 = _decodeSigs_T_11 ? 2'h0 : _decodeSigs_T_184; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_186 = _decodeSigs_T_9 ? 2'h1 : _decodeSigs_T_185; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_187 = _decodeSigs_T_7 ? 2'h1 : _decodeSigs_T_186; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_188 = _decodeSigs_T_5 ? 2'h1 : _decodeSigs_T_187; // @[Lookup.scala 34:39]
  wire [1:0] _decodeSigs_T_189 = _decodeSigs_T_3 ? 2'h1 : _decodeSigs_T_188; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_200 = _decodeSigs_T_75 ? 5'h14 : 5'h0; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_201 = _decodeSigs_T_73 ? 5'h0 : _decodeSigs_T_200; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_202 = _decodeSigs_T_71 ? 5'h0 : _decodeSigs_T_201; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_203 = _decodeSigs_T_69 ? 5'h0 : _decodeSigs_T_202; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_204 = _decodeSigs_T_67 ? 5'h0 : _decodeSigs_T_203; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_205 = _decodeSigs_T_65 ? 5'h0 : _decodeSigs_T_204; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_206 = _decodeSigs_T_63 ? 5'h0 : _decodeSigs_T_205; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_207 = _decodeSigs_T_61 ? 5'h0 : _decodeSigs_T_206; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_208 = _decodeSigs_T_59 ? 5'h0 : _decodeSigs_T_207; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_209 = _decodeSigs_T_57 ? 5'h0 : _decodeSigs_T_208; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_210 = _decodeSigs_T_55 ? 5'h0 : _decodeSigs_T_209; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_211 = _decodeSigs_T_53 ? 5'h0 : _decodeSigs_T_210; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_212 = _decodeSigs_T_51 ? 5'h0 : _decodeSigs_T_211; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_213 = _decodeSigs_T_49 ? 5'h0 : _decodeSigs_T_212; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_214 = _decodeSigs_T_47 ? 5'h0 : _decodeSigs_T_213; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_215 = _decodeSigs_T_45 ? 5'h0 : _decodeSigs_T_214; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_216 = _decodeSigs_T_43 ? 5'h0 : _decodeSigs_T_215; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_217 = _decodeSigs_T_41 ? 5'h0 : _decodeSigs_T_216; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_218 = _decodeSigs_T_39 ? 5'h0 : _decodeSigs_T_217; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_219 = _decodeSigs_T_37 ? 5'h0 : _decodeSigs_T_218; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_220 = _decodeSigs_T_35 ? 5'h8 : _decodeSigs_T_219; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_221 = _decodeSigs_T_33 ? 5'h7 : _decodeSigs_T_220; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_222 = _decodeSigs_T_31 ? 5'h6 : _decodeSigs_T_221; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_223 = _decodeSigs_T_29 ? 5'h0 : _decodeSigs_T_222; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_224 = _decodeSigs_T_27 ? 5'h0 : _decodeSigs_T_223; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_225 = _decodeSigs_T_25 ? 5'h0 : _decodeSigs_T_224; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_226 = _decodeSigs_T_23 ? 5'h0 : _decodeSigs_T_225; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_227 = _decodeSigs_T_21 ? 5'h0 : _decodeSigs_T_226; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_228 = _decodeSigs_T_19 ? 5'h0 : _decodeSigs_T_227; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_229 = _decodeSigs_T_17 ? 5'h0 : _decodeSigs_T_228; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_230 = _decodeSigs_T_15 ? 5'h0 : _decodeSigs_T_229; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_231 = _decodeSigs_T_13 ? 5'h0 : _decodeSigs_T_230; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_232 = _decodeSigs_T_11 ? 5'h0 : _decodeSigs_T_231; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_233 = _decodeSigs_T_9 ? 5'h5 : _decodeSigs_T_232; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_234 = _decodeSigs_T_7 ? 5'h4 : _decodeSigs_T_233; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_235 = _decodeSigs_T_5 ? 5'h3 : _decodeSigs_T_234; // @[Lookup.scala 34:39]
  wire [4:0] _decodeSigs_T_236 = _decodeSigs_T_3 ? 5'h2 : _decodeSigs_T_235; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_250 = _decodeSigs_T_69 ? 4'hf : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_251 = _decodeSigs_T_67 ? 4'h9 : _decodeSigs_T_250; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_252 = _decodeSigs_T_65 ? 4'h7 : _decodeSigs_T_251; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_253 = _decodeSigs_T_63 ? 4'h8 : _decodeSigs_T_252; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_254 = _decodeSigs_T_61 ? 4'h6 : _decodeSigs_T_253; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_255 = _decodeSigs_T_59 ? 4'h5 : _decodeSigs_T_254; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_256 = _decodeSigs_T_57 ? 4'he : _decodeSigs_T_255; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_257 = _decodeSigs_T_55 ? 4'h2 : _decodeSigs_T_256; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_258 = _decodeSigs_T_53 ? 4'h3 : _decodeSigs_T_257; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_259 = _decodeSigs_T_51 ? 4'hc : _decodeSigs_T_258; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_260 = _decodeSigs_T_49 ? 4'hb : _decodeSigs_T_259; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_261 = _decodeSigs_T_47 ? 4'h4 : _decodeSigs_T_260; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_262 = _decodeSigs_T_45 ? 4'h9 : _decodeSigs_T_261; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_263 = _decodeSigs_T_43 ? 4'h8 : _decodeSigs_T_262; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_264 = _decodeSigs_T_41 ? 4'ha : _decodeSigs_T_263; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_265 = _decodeSigs_T_39 ? 4'h1 : _decodeSigs_T_264; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_266 = _decodeSigs_T_37 ? 4'h0 : _decodeSigs_T_265; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_267 = _decodeSigs_T_35 ? 4'h0 : _decodeSigs_T_266; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_268 = _decodeSigs_T_33 ? 4'h0 : _decodeSigs_T_267; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_269 = _decodeSigs_T_31 ? 4'h0 : _decodeSigs_T_268; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_270 = _decodeSigs_T_29 ? 4'h0 : _decodeSigs_T_269; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_271 = _decodeSigs_T_27 ? 4'h2 : _decodeSigs_T_270; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_272 = _decodeSigs_T_25 ? 4'h3 : _decodeSigs_T_271; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_273 = _decodeSigs_T_23 ? 4'hc : _decodeSigs_T_272; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_274 = _decodeSigs_T_21 ? 4'hb : _decodeSigs_T_273; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_275 = _decodeSigs_T_19 ? 4'h4 : _decodeSigs_T_274; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_276 = _decodeSigs_T_17 ? 4'h9 : _decodeSigs_T_275; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_277 = _decodeSigs_T_15 ? 4'h8 : _decodeSigs_T_276; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_278 = _decodeSigs_T_13 ? 4'ha : _decodeSigs_T_277; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_279 = _decodeSigs_T_11 ? 4'h0 : _decodeSigs_T_278; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_280 = _decodeSigs_T_9 ? 4'h0 : _decodeSigs_T_279; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_281 = _decodeSigs_T_7 ? 4'h0 : _decodeSigs_T_280; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_282 = _decodeSigs_T_5 ? 4'h0 : _decodeSigs_T_281; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_283 = _decodeSigs_T_3 ? 4'h0 : _decodeSigs_T_282; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_284 = _decodeSigs_T_95 ? 4'h6 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_285 = _decodeSigs_T_93 ? 4'h6 : _decodeSigs_T_284; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_286 = _decodeSigs_T_91 ? 4'h6 : _decodeSigs_T_285; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_287 = _decodeSigs_T_89 ? 4'h1 : _decodeSigs_T_286; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_288 = _decodeSigs_T_87 ? 4'h1 : _decodeSigs_T_287; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_289 = _decodeSigs_T_85 ? 4'h1 : _decodeSigs_T_288; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_290 = _decodeSigs_T_83 ? 4'h0 : _decodeSigs_T_289; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_291 = _decodeSigs_T_81 ? 4'h0 : _decodeSigs_T_290; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_292 = _decodeSigs_T_79 ? 4'h0 : _decodeSigs_T_291; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_293 = _decodeSigs_T_77 ? 4'h0 : _decodeSigs_T_292; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_294 = _decodeSigs_T_75 ? 4'h0 : _decodeSigs_T_293; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_295 = _decodeSigs_T_73 ? 4'h7 : _decodeSigs_T_294; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_296 = _decodeSigs_T_71 ? 4'h1 : _decodeSigs_T_295; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_297 = _decodeSigs_T_69 ? 4'h1 : _decodeSigs_T_296; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_298 = _decodeSigs_T_67 ? 4'h1 : _decodeSigs_T_297; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_299 = _decodeSigs_T_65 ? 4'h1 : _decodeSigs_T_298; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_300 = _decodeSigs_T_63 ? 4'h1 : _decodeSigs_T_299; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_301 = _decodeSigs_T_61 ? 4'h1 : _decodeSigs_T_300; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_302 = _decodeSigs_T_59 ? 4'h1 : _decodeSigs_T_301; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_303 = _decodeSigs_T_57 ? 4'h0 : _decodeSigs_T_302; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_304 = _decodeSigs_T_55 ? 4'h1 : _decodeSigs_T_303; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_305 = _decodeSigs_T_53 ? 4'h1 : _decodeSigs_T_304; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_306 = _decodeSigs_T_51 ? 4'h1 : _decodeSigs_T_305; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_307 = _decodeSigs_T_49 ? 4'h1 : _decodeSigs_T_306; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_308 = _decodeSigs_T_47 ? 4'h1 : _decodeSigs_T_307; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_309 = _decodeSigs_T_45 ? 4'h1 : _decodeSigs_T_308; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_310 = _decodeSigs_T_43 ? 4'h1 : _decodeSigs_T_309; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_311 = _decodeSigs_T_41 ? 4'h1 : _decodeSigs_T_310; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_312 = _decodeSigs_T_39 ? 4'h1 : _decodeSigs_T_311; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_313 = _decodeSigs_T_37 ? 4'h1 : _decodeSigs_T_312; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_314 = _decodeSigs_T_35 ? 4'h1 : _decodeSigs_T_313; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_315 = _decodeSigs_T_33 ? 4'h1 : _decodeSigs_T_314; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_316 = _decodeSigs_T_31 ? 4'h1 : _decodeSigs_T_315; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_317 = _decodeSigs_T_29 ? 4'h7 : _decodeSigs_T_316; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_318 = _decodeSigs_T_27 ? 4'h1 : _decodeSigs_T_317; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_319 = _decodeSigs_T_25 ? 4'h1 : _decodeSigs_T_318; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_320 = _decodeSigs_T_23 ? 4'h1 : _decodeSigs_T_319; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_321 = _decodeSigs_T_21 ? 4'h1 : _decodeSigs_T_320; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_322 = _decodeSigs_T_19 ? 4'h1 : _decodeSigs_T_321; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_323 = _decodeSigs_T_17 ? 4'h1 : _decodeSigs_T_322; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_324 = _decodeSigs_T_15 ? 4'h1 : _decodeSigs_T_323; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_325 = _decodeSigs_T_13 ? 4'h1 : _decodeSigs_T_324; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_326 = _decodeSigs_T_11 ? 4'h1 : _decodeSigs_T_325; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_327 = _decodeSigs_T_9 ? 4'h1 : _decodeSigs_T_326; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_328 = _decodeSigs_T_7 ? 4'h1 : _decodeSigs_T_327; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_329 = _decodeSigs_T_5 ? 4'h1 : _decodeSigs_T_328; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_330 = _decodeSigs_T_3 ? 4'h1 : _decodeSigs_T_329; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_342 = _decodeSigs_T_73 ? 4'h3 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_343 = _decodeSigs_T_71 ? 4'h3 : _decodeSigs_T_342; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_344 = _decodeSigs_T_69 ? 4'h2 : _decodeSigs_T_343; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_345 = _decodeSigs_T_67 ? 4'h2 : _decodeSigs_T_344; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_346 = _decodeSigs_T_65 ? 4'h2 : _decodeSigs_T_345; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_347 = _decodeSigs_T_63 ? 4'h2 : _decodeSigs_T_346; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_348 = _decodeSigs_T_61 ? 4'h2 : _decodeSigs_T_347; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_349 = _decodeSigs_T_59 ? 4'h2 : _decodeSigs_T_348; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_350 = _decodeSigs_T_57 ? 4'h3 : _decodeSigs_T_349; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_351 = _decodeSigs_T_55 ? 4'h2 : _decodeSigs_T_350; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_352 = _decodeSigs_T_53 ? 4'h2 : _decodeSigs_T_351; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_353 = _decodeSigs_T_51 ? 4'h2 : _decodeSigs_T_352; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_354 = _decodeSigs_T_49 ? 4'h2 : _decodeSigs_T_353; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_355 = _decodeSigs_T_47 ? 4'h2 : _decodeSigs_T_354; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_356 = _decodeSigs_T_45 ? 4'h2 : _decodeSigs_T_355; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_357 = _decodeSigs_T_43 ? 4'h2 : _decodeSigs_T_356; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_358 = _decodeSigs_T_41 ? 4'h2 : _decodeSigs_T_357; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_359 = _decodeSigs_T_39 ? 4'h2 : _decodeSigs_T_358; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_360 = _decodeSigs_T_37 ? 4'h2 : _decodeSigs_T_359; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_361 = _decodeSigs_T_35 ? 4'h3 : _decodeSigs_T_360; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_362 = _decodeSigs_T_33 ? 4'h3 : _decodeSigs_T_361; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_363 = _decodeSigs_T_31 ? 4'h3 : _decodeSigs_T_362; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_364 = _decodeSigs_T_29 ? 4'h3 : _decodeSigs_T_363; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_365 = _decodeSigs_T_27 ? 4'h3 : _decodeSigs_T_364; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_366 = _decodeSigs_T_25 ? 4'h3 : _decodeSigs_T_365; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_367 = _decodeSigs_T_23 ? 4'h3 : _decodeSigs_T_366; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_368 = _decodeSigs_T_21 ? 4'h3 : _decodeSigs_T_367; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_369 = _decodeSigs_T_19 ? 4'h3 : _decodeSigs_T_368; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_370 = _decodeSigs_T_17 ? 4'h3 : _decodeSigs_T_369; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_371 = _decodeSigs_T_15 ? 4'h3 : _decodeSigs_T_370; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_372 = _decodeSigs_T_13 ? 4'h3 : _decodeSigs_T_371; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_373 = _decodeSigs_T_11 ? 4'h3 : _decodeSigs_T_372; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_374 = _decodeSigs_T_9 ? 4'h3 : _decodeSigs_T_373; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_375 = _decodeSigs_T_7 ? 4'h3 : _decodeSigs_T_374; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_376 = _decodeSigs_T_5 ? 4'h3 : _decodeSigs_T_375; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_377 = _decodeSigs_T_3 ? 4'h3 : _decodeSigs_T_376; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_378 = _decodeSigs_T_95 ? 3'h5 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_379 = _decodeSigs_T_93 ? 3'h5 : _decodeSigs_T_378; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_380 = _decodeSigs_T_91 ? 3'h5 : _decodeSigs_T_379; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_381 = _decodeSigs_T_89 ? 3'h0 : _decodeSigs_T_380; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_382 = _decodeSigs_T_87 ? 3'h0 : _decodeSigs_T_381; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_383 = _decodeSigs_T_85 ? 3'h0 : _decodeSigs_T_382; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_384 = _decodeSigs_T_83 ? 3'h0 : _decodeSigs_T_383; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_385 = _decodeSigs_T_81 ? 3'h0 : _decodeSigs_T_384; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_386 = _decodeSigs_T_79 ? 3'h0 : _decodeSigs_T_385; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_387 = _decodeSigs_T_77 ? 3'h0 : _decodeSigs_T_386; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_388 = _decodeSigs_T_75 ? 3'h0 : _decodeSigs_T_387; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_389 = _decodeSigs_T_73 ? 3'h4 : _decodeSigs_T_388; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_390 = _decodeSigs_T_71 ? 3'h0 : _decodeSigs_T_389; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_391 = _decodeSigs_T_69 ? 3'h2 : _decodeSigs_T_390; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_392 = _decodeSigs_T_67 ? 3'h2 : _decodeSigs_T_391; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_393 = _decodeSigs_T_65 ? 3'h2 : _decodeSigs_T_392; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_394 = _decodeSigs_T_63 ? 3'h2 : _decodeSigs_T_393; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_395 = _decodeSigs_T_61 ? 3'h2 : _decodeSigs_T_394; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_396 = _decodeSigs_T_59 ? 3'h2 : _decodeSigs_T_395; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_397 = _decodeSigs_T_57 ? 3'h3 : _decodeSigs_T_396; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_398 = _decodeSigs_T_55 ? 3'h0 : _decodeSigs_T_397; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_399 = _decodeSigs_T_53 ? 3'h0 : _decodeSigs_T_398; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_400 = _decodeSigs_T_51 ? 3'h0 : _decodeSigs_T_399; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_401 = _decodeSigs_T_49 ? 3'h0 : _decodeSigs_T_400; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_402 = _decodeSigs_T_47 ? 3'h0 : _decodeSigs_T_401; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_403 = _decodeSigs_T_45 ? 3'h0 : _decodeSigs_T_402; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_404 = _decodeSigs_T_43 ? 3'h0 : _decodeSigs_T_403; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_405 = _decodeSigs_T_41 ? 3'h0 : _decodeSigs_T_404; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_406 = _decodeSigs_T_39 ? 3'h0 : _decodeSigs_T_405; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_407 = _decodeSigs_T_37 ? 3'h0 : _decodeSigs_T_406; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_408 = _decodeSigs_T_35 ? 3'h1 : _decodeSigs_T_407; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_409 = _decodeSigs_T_33 ? 3'h1 : _decodeSigs_T_408; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_410 = _decodeSigs_T_31 ? 3'h1 : _decodeSigs_T_409; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_411 = _decodeSigs_T_29 ? 3'h3 : _decodeSigs_T_410; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_412 = _decodeSigs_T_27 ? 3'h0 : _decodeSigs_T_411; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_413 = _decodeSigs_T_25 ? 3'h0 : _decodeSigs_T_412; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_414 = _decodeSigs_T_23 ? 3'h0 : _decodeSigs_T_413; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_415 = _decodeSigs_T_21 ? 3'h0 : _decodeSigs_T_414; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_416 = _decodeSigs_T_19 ? 3'h0 : _decodeSigs_T_415; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_417 = _decodeSigs_T_17 ? 3'h0 : _decodeSigs_T_416; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_418 = _decodeSigs_T_15 ? 3'h0 : _decodeSigs_T_417; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_419 = _decodeSigs_T_13 ? 3'h0 : _decodeSigs_T_418; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_420 = _decodeSigs_T_11 ? 3'h0 : _decodeSigs_T_419; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_421 = _decodeSigs_T_9 ? 3'h0 : _decodeSigs_T_420; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_422 = _decodeSigs_T_7 ? 3'h0 : _decodeSigs_T_421; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_423 = _decodeSigs_T_5 ? 3'h0 : _decodeSigs_T_422; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_424 = _decodeSigs_T_3 ? 3'h0 : _decodeSigs_T_423; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_425 = _decodeSigs_T_95 ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_426 = _decodeSigs_T_93 ? 1'h0 : _decodeSigs_T_425; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_427 = _decodeSigs_T_91 ? 1'h0 : _decodeSigs_T_426; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_428 = _decodeSigs_T_89 ? 1'h0 : _decodeSigs_T_427; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_429 = _decodeSigs_T_87 ? 1'h0 : _decodeSigs_T_428; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_430 = _decodeSigs_T_85 ? 1'h0 : _decodeSigs_T_429; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_431 = _decodeSigs_T_83 ? 1'h0 : _decodeSigs_T_430; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_432 = _decodeSigs_T_81 ? 1'h0 : _decodeSigs_T_431; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_433 = _decodeSigs_T_79 ? 1'h0 : _decodeSigs_T_432; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_434 = _decodeSigs_T_77 ? 1'h0 : _decodeSigs_T_433; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_444 = _decodeSigs_T_57 ? 1'h0 : _decodeSigs_T_59 | (_decodeSigs_T_61 | (_decodeSigs_T_63 | (
    _decodeSigs_T_65 | (_decodeSigs_T_67 | (_decodeSigs_T_69 | (_decodeSigs_T_71 | (_decodeSigs_T_73 | (_decodeSigs_T_75
     | _decodeSigs_T_434)))))))); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_445 = _decodeSigs_T_55 ? 1'h0 : _decodeSigs_T_444; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_446 = _decodeSigs_T_53 ? 1'h0 : _decodeSigs_T_445; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_447 = _decodeSigs_T_51 ? 1'h0 : _decodeSigs_T_446; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_448 = _decodeSigs_T_49 ? 1'h0 : _decodeSigs_T_447; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_449 = _decodeSigs_T_47 ? 1'h0 : _decodeSigs_T_448; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_450 = _decodeSigs_T_45 ? 1'h0 : _decodeSigs_T_449; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_451 = _decodeSigs_T_43 ? 1'h0 : _decodeSigs_T_450; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_452 = _decodeSigs_T_41 ? 1'h0 : _decodeSigs_T_451; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_453 = _decodeSigs_T_39 ? 1'h0 : _decodeSigs_T_452; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_454 = _decodeSigs_T_37 ? 1'h0 : _decodeSigs_T_453; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_458 = _decodeSigs_T_29 ? 1'h0 : _decodeSigs_T_31 | (_decodeSigs_T_33 | (_decodeSigs_T_35 |
    _decodeSigs_T_454)); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_462 = _decodeSigs_T_21 ? 1'h0 : _decodeSigs_T_23 | (_decodeSigs_T_25 | (_decodeSigs_T_27 |
    _decodeSigs_T_458)); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_466 = _decodeSigs_T_13 ? 1'h0 : _decodeSigs_T_15 | (_decodeSigs_T_17 | (_decodeSigs_T_19 |
    _decodeSigs_T_462)); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_478 = _decodeSigs_T_83 ? 1'h0 : _decodeSigs_T_85 | (_decodeSigs_T_87 | (_decodeSigs_T_89 | (
    _decodeSigs_T_91 | (_decodeSigs_T_93 | _decodeSigs_T_95)))); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_479 = _decodeSigs_T_81 ? 1'h0 : _decodeSigs_T_478; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_480 = _decodeSigs_T_79 ? 1'h0 : _decodeSigs_T_479; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_481 = _decodeSigs_T_77 ? 1'h0 : _decodeSigs_T_480; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_482 = _decodeSigs_T_75 ? 1'h0 : _decodeSigs_T_481; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_485 = _decodeSigs_T_69 ? 1'h0 : _decodeSigs_T_71 | (_decodeSigs_T_73 | _decodeSigs_T_482); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_486 = _decodeSigs_T_67 ? 1'h0 : _decodeSigs_T_485; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_487 = _decodeSigs_T_65 ? 1'h0 : _decodeSigs_T_486; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_488 = _decodeSigs_T_63 ? 1'h0 : _decodeSigs_T_487; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_489 = _decodeSigs_T_61 ? 1'h0 : _decodeSigs_T_488; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_490 = _decodeSigs_T_59 ? 1'h0 : _decodeSigs_T_489; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_502 = _decodeSigs_T_35 ? 1'h0 : _decodeSigs_T_37 | (_decodeSigs_T_39 | (_decodeSigs_T_41 | (
    _decodeSigs_T_43 | (_decodeSigs_T_45 | (_decodeSigs_T_47 | (_decodeSigs_T_49 | (_decodeSigs_T_51 | (_decodeSigs_T_53
     | (_decodeSigs_T_55 | (_decodeSigs_T_57 | _decodeSigs_T_490)))))))))); // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_503 = _decodeSigs_T_33 ? 1'h0 : _decodeSigs_T_502; // @[Lookup.scala 34:39]
  wire  _decodeSigs_T_504 = _decodeSigs_T_31 ? 1'h0 : _decodeSigs_T_503; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_520 = _decodeSigs_T_93 ? 3'h4 : _decodeSigs_T_378; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_521 = _decodeSigs_T_91 ? 3'h3 : _decodeSigs_T_520; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_522 = _decodeSigs_T_89 ? 3'h5 : _decodeSigs_T_521; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_523 = _decodeSigs_T_87 ? 3'h4 : _decodeSigs_T_522; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_524 = _decodeSigs_T_85 ? 3'h3 : _decodeSigs_T_523; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_525 = _decodeSigs_T_83 ? 3'h0 : _decodeSigs_T_524; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_526 = _decodeSigs_T_81 ? 3'h0 : _decodeSigs_T_525; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_527 = _decodeSigs_T_79 ? 3'h0 : _decodeSigs_T_526; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_528 = _decodeSigs_T_77 ? 3'h0 : _decodeSigs_T_527; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_529 = _decodeSigs_T_75 ? 3'h0 : _decodeSigs_T_528; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_530 = _decodeSigs_T_73 ? 3'h0 : _decodeSigs_T_529; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_531 = _decodeSigs_T_71 ? 3'h0 : _decodeSigs_T_530; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_532 = _decodeSigs_T_69 ? 3'h0 : _decodeSigs_T_531; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_533 = _decodeSigs_T_67 ? 3'h0 : _decodeSigs_T_532; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_534 = _decodeSigs_T_65 ? 3'h0 : _decodeSigs_T_533; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_535 = _decodeSigs_T_63 ? 3'h0 : _decodeSigs_T_534; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_536 = _decodeSigs_T_61 ? 3'h0 : _decodeSigs_T_535; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_537 = _decodeSigs_T_59 ? 3'h0 : _decodeSigs_T_536; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_538 = _decodeSigs_T_57 ? 3'h0 : _decodeSigs_T_537; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_539 = _decodeSigs_T_55 ? 3'h0 : _decodeSigs_T_538; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_540 = _decodeSigs_T_53 ? 3'h0 : _decodeSigs_T_539; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_541 = _decodeSigs_T_51 ? 3'h0 : _decodeSigs_T_540; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_542 = _decodeSigs_T_49 ? 3'h0 : _decodeSigs_T_541; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_543 = _decodeSigs_T_47 ? 3'h0 : _decodeSigs_T_542; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_544 = _decodeSigs_T_45 ? 3'h0 : _decodeSigs_T_543; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_545 = _decodeSigs_T_43 ? 3'h0 : _decodeSigs_T_544; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_546 = _decodeSigs_T_41 ? 3'h0 : _decodeSigs_T_545; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_547 = _decodeSigs_T_39 ? 3'h0 : _decodeSigs_T_546; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_548 = _decodeSigs_T_37 ? 3'h0 : _decodeSigs_T_547; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_549 = _decodeSigs_T_35 ? 3'h0 : _decodeSigs_T_548; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_550 = _decodeSigs_T_33 ? 3'h0 : _decodeSigs_T_549; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_551 = _decodeSigs_T_31 ? 3'h0 : _decodeSigs_T_550; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_552 = _decodeSigs_T_29 ? 3'h0 : _decodeSigs_T_551; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_553 = _decodeSigs_T_27 ? 3'h0 : _decodeSigs_T_552; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_554 = _decodeSigs_T_25 ? 3'h0 : _decodeSigs_T_553; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_555 = _decodeSigs_T_23 ? 3'h0 : _decodeSigs_T_554; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_556 = _decodeSigs_T_21 ? 3'h0 : _decodeSigs_T_555; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_557 = _decodeSigs_T_19 ? 3'h0 : _decodeSigs_T_556; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_558 = _decodeSigs_T_17 ? 3'h0 : _decodeSigs_T_557; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_559 = _decodeSigs_T_15 ? 3'h0 : _decodeSigs_T_558; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_560 = _decodeSigs_T_13 ? 3'h0 : _decodeSigs_T_559; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_561 = _decodeSigs_T_11 ? 3'h0 : _decodeSigs_T_560; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_562 = _decodeSigs_T_9 ? 3'h0 : _decodeSigs_T_561; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_563 = _decodeSigs_T_7 ? 3'h0 : _decodeSigs_T_562; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_564 = _decodeSigs_T_5 ? 3'h0 : _decodeSigs_T_563; // @[Lookup.scala 34:39]
  wire [2:0] _decodeSigs_T_565 = _decodeSigs_T_3 ? 3'h0 : _decodeSigs_T_564; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_566 = _decodeSigs_T_95 ? 4'h0 : 4'h5; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_567 = _decodeSigs_T_93 ? 4'h0 : _decodeSigs_T_566; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_568 = _decodeSigs_T_91 ? 4'h0 : _decodeSigs_T_567; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_569 = _decodeSigs_T_89 ? 4'h0 : _decodeSigs_T_568; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_570 = _decodeSigs_T_87 ? 4'h0 : _decodeSigs_T_569; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_571 = _decodeSigs_T_85 ? 4'h0 : _decodeSigs_T_570; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_572 = _decodeSigs_T_83 ? 4'h3 : _decodeSigs_T_571; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_573 = _decodeSigs_T_81 ? 4'h4 : _decodeSigs_T_572; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_574 = _decodeSigs_T_79 ? 4'h2 : _decodeSigs_T_573; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_575 = _decodeSigs_T_77 ? 4'h1 : _decodeSigs_T_574; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_576 = _decodeSigs_T_75 ? 4'h0 : _decodeSigs_T_575; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_577 = _decodeSigs_T_73 ? 4'h0 : _decodeSigs_T_576; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_578 = _decodeSigs_T_71 ? 4'h0 : _decodeSigs_T_577; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_579 = _decodeSigs_T_69 ? 4'h0 : _decodeSigs_T_578; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_580 = _decodeSigs_T_67 ? 4'h0 : _decodeSigs_T_579; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_581 = _decodeSigs_T_65 ? 4'h0 : _decodeSigs_T_580; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_582 = _decodeSigs_T_63 ? 4'h0 : _decodeSigs_T_581; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_583 = _decodeSigs_T_61 ? 4'h0 : _decodeSigs_T_582; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_584 = _decodeSigs_T_59 ? 4'h0 : _decodeSigs_T_583; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_585 = _decodeSigs_T_57 ? 4'h0 : _decodeSigs_T_584; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_586 = _decodeSigs_T_55 ? 4'h0 : _decodeSigs_T_585; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_587 = _decodeSigs_T_53 ? 4'h0 : _decodeSigs_T_586; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_588 = _decodeSigs_T_51 ? 4'h0 : _decodeSigs_T_587; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_589 = _decodeSigs_T_49 ? 4'h0 : _decodeSigs_T_588; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_590 = _decodeSigs_T_47 ? 4'h0 : _decodeSigs_T_589; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_591 = _decodeSigs_T_45 ? 4'h0 : _decodeSigs_T_590; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_592 = _decodeSigs_T_43 ? 4'h0 : _decodeSigs_T_591; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_593 = _decodeSigs_T_41 ? 4'h0 : _decodeSigs_T_592; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_594 = _decodeSigs_T_39 ? 4'h0 : _decodeSigs_T_593; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_595 = _decodeSigs_T_37 ? 4'h0 : _decodeSigs_T_594; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_596 = _decodeSigs_T_35 ? 4'h0 : _decodeSigs_T_595; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_597 = _decodeSigs_T_33 ? 4'h0 : _decodeSigs_T_596; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_598 = _decodeSigs_T_31 ? 4'h0 : _decodeSigs_T_597; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_599 = _decodeSigs_T_29 ? 4'h0 : _decodeSigs_T_598; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_600 = _decodeSigs_T_27 ? 4'h0 : _decodeSigs_T_599; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_601 = _decodeSigs_T_25 ? 4'h0 : _decodeSigs_T_600; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_602 = _decodeSigs_T_23 ? 4'h0 : _decodeSigs_T_601; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_603 = _decodeSigs_T_21 ? 4'h0 : _decodeSigs_T_602; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_604 = _decodeSigs_T_19 ? 4'h0 : _decodeSigs_T_603; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_605 = _decodeSigs_T_17 ? 4'h0 : _decodeSigs_T_604; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_606 = _decodeSigs_T_15 ? 4'h0 : _decodeSigs_T_605; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_607 = _decodeSigs_T_13 ? 4'h0 : _decodeSigs_T_606; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_608 = _decodeSigs_T_11 ? 4'h0 : _decodeSigs_T_607; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_609 = _decodeSigs_T_9 ? 4'h0 : _decodeSigs_T_608; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_610 = _decodeSigs_T_7 ? 4'h0 : _decodeSigs_T_609; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_611 = _decodeSigs_T_5 ? 4'h0 : _decodeSigs_T_610; // @[Lookup.scala 34:39]
  wire [3:0] _decodeSigs_T_612 = _decodeSigs_T_3 ? 4'h0 : _decodeSigs_T_611; // @[Lookup.scala 34:39]
  assign io_out_isBranch = _decodeSigs_T_1 ? 1'h0 : _decodeSigs_T_142; // @[Lookup.scala 34:39]
  assign io_out_resultSrc = _decodeSigs_T_1 ? 2'h1 : _decodeSigs_T_189; // @[Lookup.scala 34:39]
  assign io_out_aluOpSel = _decodeSigs_T_1 ? 4'h0 : _decodeSigs_T_283; // @[Lookup.scala 34:39]
  assign io_out_lsuOp = _decodeSigs_T_1 ? 5'h1 : _decodeSigs_T_236; // @[Lookup.scala 34:39]
  assign io_out_aluSrc1 = _decodeSigs_T_1 ? 4'h1 : _decodeSigs_T_330; // @[Lookup.scala 34:39]
  assign io_out_aluSrc2 = _decodeSigs_T_1 ? 4'h3 : _decodeSigs_T_377; // @[Lookup.scala 34:39]
  assign io_out_immSrc = _decodeSigs_T_1 ? 3'h0 : _decodeSigs_T_424; // @[Lookup.scala 34:39]
  assign io_out_immSign = _decodeSigs_T_1 | (_decodeSigs_T_3 | (_decodeSigs_T_5 | (_decodeSigs_T_7 | (_decodeSigs_T_9 |
    (_decodeSigs_T_11 | _decodeSigs_T_466))))); // @[Lookup.scala 34:39]
  assign io_out_regWrEn = _decodeSigs_T_1 | (_decodeSigs_T_3 | (_decodeSigs_T_5 | (_decodeSigs_T_7 | (_decodeSigs_T_9 |
    (_decodeSigs_T_11 | (_decodeSigs_T_13 | (_decodeSigs_T_15 | (_decodeSigs_T_17 | (_decodeSigs_T_19 | (
    _decodeSigs_T_21 | (_decodeSigs_T_23 | (_decodeSigs_T_25 | (_decodeSigs_T_27 | (_decodeSigs_T_29 | _decodeSigs_T_504
    )))))))))))))); // @[Lookup.scala 34:39]
  assign io_out_csrOp = _decodeSigs_T_1 ? 3'h0 : _decodeSigs_T_565; // @[Lookup.scala 34:39]
  assign io_out_excType = _decodeSigs_T_1 ? 4'h0 : _decodeSigs_T_612; // @[Lookup.scala 34:39]
endmodule
module CtrlUnit(
  output        io_out_isBranch,
  output        io_out_isJump,
  output [1:0]  io_out_resultSrc,
  output [3:0]  io_out_aluOpSel,
  output [4:0]  io_out_lsuOp,
  output [3:0]  io_out_aluSrc1,
  output [3:0]  io_out_aluSrc2,
  output [2:0]  io_out_immSrc,
  output        io_out_immSign,
  output        io_out_regWrEn,
  output        io_out_pcAddReg,
  output [2:0]  io_out_csrOp,
  output [3:0]  io_out_excType,
  input  [31:0] io_in_inst
);
  wire [31:0] decoder_io_inst; // @[CtrlUnit.scala 59:25]
  wire  decoder_io_out_isBranch; // @[CtrlUnit.scala 59:25]
  wire [1:0] decoder_io_out_resultSrc; // @[CtrlUnit.scala 59:25]
  wire [3:0] decoder_io_out_aluOpSel; // @[CtrlUnit.scala 59:25]
  wire [4:0] decoder_io_out_lsuOp; // @[CtrlUnit.scala 59:25]
  wire [3:0] decoder_io_out_aluSrc1; // @[CtrlUnit.scala 59:25]
  wire [3:0] decoder_io_out_aluSrc2; // @[CtrlUnit.scala 59:25]
  wire [2:0] decoder_io_out_immSrc; // @[CtrlUnit.scala 59:25]
  wire  decoder_io_out_immSign; // @[CtrlUnit.scala 59:25]
  wire  decoder_io_out_regWrEn; // @[CtrlUnit.scala 59:25]
  wire [2:0] decoder_io_out_csrOp; // @[CtrlUnit.scala 59:25]
  wire [3:0] decoder_io_out_excType; // @[CtrlUnit.scala 59:25]
  wire [6:0] opcode = io_in_inst[6:0]; // @[util.scala 74:34]
  wire  _io_out_pcAddReg_T_1 = 7'h67 == opcode; // @[CtrlUnit.scala 81:31]
  Decoder decoder ( // @[CtrlUnit.scala 59:25]
    .io_inst(decoder_io_inst),
    .io_out_isBranch(decoder_io_out_isBranch),
    .io_out_resultSrc(decoder_io_out_resultSrc),
    .io_out_aluOpSel(decoder_io_out_aluOpSel),
    .io_out_lsuOp(decoder_io_out_lsuOp),
    .io_out_aluSrc1(decoder_io_out_aluSrc1),
    .io_out_aluSrc2(decoder_io_out_aluSrc2),
    .io_out_immSrc(decoder_io_out_immSrc),
    .io_out_immSign(decoder_io_out_immSign),
    .io_out_regWrEn(decoder_io_out_regWrEn),
    .io_out_csrOp(decoder_io_out_csrOp),
    .io_out_excType(decoder_io_out_excType)
  );
  assign io_out_isBranch = decoder_io_out_isBranch; // @[CtrlUnit.scala 63:21]
  assign io_out_isJump = _io_out_pcAddReg_T_1 | 7'h6f == opcode; // @[CtrlUnit.scala 82:45]
  assign io_out_resultSrc = decoder_io_out_resultSrc; // @[CtrlUnit.scala 64:21]
  assign io_out_aluOpSel = decoder_io_out_aluOpSel; // @[CtrlUnit.scala 67:21]
  assign io_out_lsuOp = decoder_io_out_lsuOp; // @[CtrlUnit.scala 68:21]
  assign io_out_aluSrc1 = decoder_io_out_aluSrc1; // @[CtrlUnit.scala 70:21]
  assign io_out_aluSrc2 = decoder_io_out_aluSrc2; // @[CtrlUnit.scala 71:21]
  assign io_out_immSrc = decoder_io_out_immSrc; // @[CtrlUnit.scala 72:21]
  assign io_out_immSign = decoder_io_out_immSign; // @[CtrlUnit.scala 73:21]
  assign io_out_regWrEn = decoder_io_out_regWrEn; // @[CtrlUnit.scala 74:21]
  assign io_out_pcAddReg = 7'h67 == opcode; // @[CtrlUnit.scala 81:31]
  assign io_out_csrOp = decoder_io_out_csrOp; // @[CtrlUnit.scala 76:21]
  assign io_out_excType = decoder_io_out_excType; // @[CtrlUnit.scala 77:21]
  assign decoder_io_inst = io_in_inst; // @[CtrlUnit.scala 61:27]
endmodule
module ImmGen(
  input  [31:0] io_inst,
  input  [2:0]  io_immSrc,
  input         io_immSign,
  output [31:0] io_imm
);
  wire [31:0] immI = {{20'd0}, io_inst[31:20]}; // @[util.scala 62:36]
  wire [11:0] _immS_T_2 = {io_inst[31:25],io_inst[11:7]}; // @[Cat.scala 33:92]
  wire [31:0] immS = {{20'd0}, _immS_T_2}; // @[util.scala 62:36]
  wire [12:0] _immB_T_4 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] immB = {{19'd0}, _immB_T_4}; // @[util.scala 62:36]
  wire [31:0] immU = {io_inst[31:12], 12'h0}; // @[ImmGen.scala 26:36]
  wire [20:0] _immJ_T_4 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] immJ = {{11'd0}, _immJ_T_4}; // @[util.scala 62:36]
  wire [11:0] _immI_S_T_1 = io_inst[31:20]; // @[util.scala 51:20]
  wire  immI_S_signBit = _immI_S_T_1[11]; // @[util.scala 42:27]
  wire [9:0] immI_S_out_lo = {immI_S_signBit,immI_S_signBit,immI_S_signBit,immI_S_signBit,immI_S_signBit,immI_S_signBit,
    immI_S_signBit,immI_S_signBit,immI_S_signBit,immI_S_signBit}; // @[Cat.scala 33:92]
  wire [11:0] _immI_S_out_T_1 = io_inst[31:20]; // @[util.scala 46:75]
  wire [31:0] immI_S = {immI_S_out_lo,immI_S_out_lo,_immI_S_out_T_1}; // @[Cat.scala 33:92]
  wire [11:0] _immS_S_T_3 = {io_inst[31:25],io_inst[11:7]}; // @[util.scala 51:20]
  wire  immS_S_signBit = _immS_S_T_3[11]; // @[util.scala 42:27]
  wire [9:0] immS_S_out_lo = {immS_S_signBit,immS_S_signBit,immS_S_signBit,immS_S_signBit,immS_S_signBit,immS_S_signBit,
    immS_S_signBit,immS_S_signBit,immS_S_signBit,immS_S_signBit}; // @[Cat.scala 33:92]
  wire [11:0] _immS_S_out_T_1 = {io_inst[31:25],io_inst[11:7]}; // @[util.scala 46:75]
  wire [31:0] immS_S = {immS_S_out_lo,immS_S_out_lo,_immS_S_out_T_1}; // @[Cat.scala 33:92]
  wire [12:0] _immB_S_T_5 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[util.scala 51:20]
  wire  immB_S_signBit = _immB_S_T_5[12]; // @[util.scala 42:27]
  wire [9:0] immB_S_out_hi = {immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,
    immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit}; // @[Cat.scala 33:92]
  wire [18:0] _immB_S_out_T = {immB_S_out_hi,immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit,
    immB_S_signBit,immB_S_signBit,immB_S_signBit,immB_S_signBit}; // @[Cat.scala 33:92]
  wire [12:0] _immB_S_out_T_1 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[util.scala 46:75]
  wire [31:0] immB_S = {_immB_S_out_T,_immB_S_out_T_1}; // @[Cat.scala 33:92]
  wire [31:0] immU_S = {io_inst[31:12], 12'h0}; // @[util.scala 44:18]
  wire [20:0] _immJ_S_T_5 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[util.scala 51:20]
  wire  immJ_S_signBit = _immJ_S_T_5[20]; // @[util.scala 42:27]
  wire [4:0] immJ_S_out_lo = {immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit}; // @[Cat.scala 33:92]
  wire [20:0] _immJ_S_out_T_1 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[util.scala 46:75]
  wire [31:0] immJ_S = {immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,immJ_S_signBit,
    immJ_S_out_lo,_immJ_S_out_T_1}; // @[Cat.scala 33:92]
  wire [31:0] _out_T_3 = 3'h1 == io_immSrc ? immS_S : immI_S; // @[Mux.scala 81:58]
  wire [31:0] _out_T_5 = 3'h2 == io_immSrc ? immB_S : _out_T_3; // @[Mux.scala 81:58]
  wire [31:0] _out_T_7 = 3'h3 == io_immSrc ? immU_S : _out_T_5; // @[Mux.scala 81:58]
  wire [31:0] _out_T_9 = 3'h4 == io_immSrc ? immJ_S : _out_T_7; // @[Mux.scala 81:58]
  wire [31:0] _out_T_13 = 3'h1 == io_immSrc ? immS : immI; // @[Mux.scala 81:58]
  wire [31:0] _out_T_15 = 3'h2 == io_immSrc ? immB : _out_T_13; // @[Mux.scala 81:58]
  wire [31:0] _out_T_17 = 3'h3 == io_immSrc ? immU : _out_T_15; // @[Mux.scala 81:58]
  wire [31:0] _out_T_19 = 3'h4 == io_immSrc ? immJ : _out_T_17; // @[Mux.scala 81:58]
  wire [31:0] _GEN_0 = io_immSign ? _out_T_9 : _out_T_19; // @[ImmGen.scala 37:19 38:13 46:13]
  wire [31:0] out_out = {{27'd0}, io_inst[19:15]}; // @[util.scala 62:36]
  assign io_imm = io_immSrc == 3'h5 ? out_out : _GEN_0; // @[ImmGen.scala 55:30 56:13]
endmodule
module Decode(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_pcNext4,
  input         io_in_bits_instState_commit,
  input  [31:0] io_in_bits_instState_pc,
  input  [31:0] io_in_bits_instState_inst,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_isBranch,
  output        io_out_bits_isJump,
  output [1:0]  io_out_bits_resultSrc,
  output [4:0]  io_out_bits_lsuOp,
  output [3:0]  io_out_bits_aluOpSel,
  output        io_out_bits_immSign,
  output        io_out_bits_regWrEn,
  output        io_out_bits_pcAddReg,
  output [31:0] io_out_bits_pcNext4,
  output [31:0] io_out_bits_aluIn1,
  output [31:0] io_out_bits_aluIn2,
  output        io_out_bits_aluIn1IsReg,
  output        io_out_bits_aluIn2IsReg,
  output [31:0] io_out_bits_imm,
  output [31:0] io_out_bits_data2,
  output [3:0]  io_out_bits_excType,
  output [2:0]  io_out_bits_csrOp,
  output        io_out_bits_instState_commit,
  output [31:0] io_out_bits_instState_pc,
  output [31:0] io_out_bits_instState_inst,
  output [4:0]  io_hazard_out_rs1,
  output [4:0]  io_hazard_out_rs2,
  input         io_hazard_in_stall,
  output [4:0]  io_regfile_rs1,
  output [4:0]  io_regfile_rs2,
  input  [31:0] io_regfile_rdata1,
  input  [31:0] io_regfile_rdata2,
  input         io_ctrl_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ctrlUnit_io_out_isBranch; // @[2_Decode.scala 119:29]
  wire  ctrlUnit_io_out_isJump; // @[2_Decode.scala 119:29]
  wire [1:0] ctrlUnit_io_out_resultSrc; // @[2_Decode.scala 119:29]
  wire [3:0] ctrlUnit_io_out_aluOpSel; // @[2_Decode.scala 119:29]
  wire [4:0] ctrlUnit_io_out_lsuOp; // @[2_Decode.scala 119:29]
  wire [3:0] ctrlUnit_io_out_aluSrc1; // @[2_Decode.scala 119:29]
  wire [3:0] ctrlUnit_io_out_aluSrc2; // @[2_Decode.scala 119:29]
  wire [2:0] ctrlUnit_io_out_immSrc; // @[2_Decode.scala 119:29]
  wire  ctrlUnit_io_out_immSign; // @[2_Decode.scala 119:29]
  wire  ctrlUnit_io_out_regWrEn; // @[2_Decode.scala 119:29]
  wire  ctrlUnit_io_out_pcAddReg; // @[2_Decode.scala 119:29]
  wire [2:0] ctrlUnit_io_out_csrOp; // @[2_Decode.scala 119:29]
  wire [3:0] ctrlUnit_io_out_excType; // @[2_Decode.scala 119:29]
  wire [31:0] ctrlUnit_io_in_inst; // @[2_Decode.scala 119:29]
  wire [31:0] immGen_io_inst; // @[2_Decode.scala 142:24]
  wire [2:0] immGen_io_immSrc; // @[2_Decode.scala 142:24]
  wire  immGen_io_immSign; // @[2_Decode.scala 142:24]
  wire [31:0] immGen_io_imm; // @[2_Decode.scala 142:24]
  wire  _io_in_ready_T = ~io_hazard_in_stall; // @[2_Decode.scala 79:20]
  wire  _io_in_ready_T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire  decodeLatch = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  reg [31:0] stageReg_pcNext4; // @[2_Decode.scala 82:27]
  reg  stageReg_instState_commit; // @[2_Decode.scala 82:27]
  reg [31:0] stageReg_instState_pc; // @[2_Decode.scala 82:27]
  reg [31:0] stageReg_instState_inst; // @[2_Decode.scala 82:27]
  wire [4:0] rs1 = stageReg_instState_inst[19:15]; // @[util.scala 72:31]
  wire [31:0] io_out_bits_aluIn1_out = {{27'd0}, rs1}; // @[util.scala 62:36]
  wire [31:0] _io_out_bits_aluIn1_T_1 = 4'h1 == ctrlUnit_io_out_aluSrc1 ? io_regfile_rdata1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_bits_aluIn1_T_3 = 4'h2 == ctrlUnit_io_out_aluSrc1 ? io_regfile_rdata2 : _io_out_bits_aluIn1_T_1; // @[Mux.scala 81:58]
  wire [31:0] imm = immGen_io_imm; // @[2_Decode.scala 146:25 96:25]
  wire [31:0] _io_out_bits_aluIn1_T_5 = 4'h3 == ctrlUnit_io_out_aluSrc1 ? imm : _io_out_bits_aluIn1_T_3; // @[Mux.scala 81:58]
  wire [31:0] _io_out_bits_aluIn1_T_7 = 4'h6 == ctrlUnit_io_out_aluSrc1 ? io_out_bits_aluIn1_out :
    _io_out_bits_aluIn1_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_out_bits_aluIn1_T_9 = 4'h7 == ctrlUnit_io_out_aluSrc1 ? stageReg_instState_pc :
    _io_out_bits_aluIn1_T_7; // @[Mux.scala 81:58]
  wire [31:0] _io_out_bits_aluIn2_T_1 = 4'h1 == ctrlUnit_io_out_aluSrc2 ? io_regfile_rdata1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_bits_aluIn2_T_3 = 4'h2 == ctrlUnit_io_out_aluSrc2 ? io_regfile_rdata2 : _io_out_bits_aluIn2_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_out_bits_aluIn2_T_5 = 4'h3 == ctrlUnit_io_out_aluSrc2 ? imm : _io_out_bits_aluIn2_T_3; // @[Mux.scala 81:58]
  wire [31:0] _io_out_bits_aluIn2_T_7 = 4'h6 == ctrlUnit_io_out_aluSrc2 ? io_out_bits_aluIn1_out :
    _io_out_bits_aluIn2_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_out_bits_aluIn2_T_9 = 4'h7 == ctrlUnit_io_out_aluSrc2 ? stageReg_instState_pc :
    _io_out_bits_aluIn2_T_7; // @[Mux.scala 81:58]
  CtrlUnit ctrlUnit ( // @[2_Decode.scala 119:29]
    .io_out_isBranch(ctrlUnit_io_out_isBranch),
    .io_out_isJump(ctrlUnit_io_out_isJump),
    .io_out_resultSrc(ctrlUnit_io_out_resultSrc),
    .io_out_aluOpSel(ctrlUnit_io_out_aluOpSel),
    .io_out_lsuOp(ctrlUnit_io_out_lsuOp),
    .io_out_aluSrc1(ctrlUnit_io_out_aluSrc1),
    .io_out_aluSrc2(ctrlUnit_io_out_aluSrc2),
    .io_out_immSrc(ctrlUnit_io_out_immSrc),
    .io_out_immSign(ctrlUnit_io_out_immSign),
    .io_out_regWrEn(ctrlUnit_io_out_regWrEn),
    .io_out_pcAddReg(ctrlUnit_io_out_pcAddReg),
    .io_out_csrOp(ctrlUnit_io_out_csrOp),
    .io_out_excType(ctrlUnit_io_out_excType),
    .io_in_inst(ctrlUnit_io_in_inst)
  );
  ImmGen immGen ( // @[2_Decode.scala 142:24]
    .io_inst(immGen_io_inst),
    .io_immSrc(immGen_io_immSrc),
    .io_immSign(immGen_io_immSign),
    .io_imm(immGen_io_imm)
  );
  assign io_in_ready = ~io_hazard_in_stall & io_in_valid & _io_in_ready_T_2; // @[2_Decode.scala 79:42]
  assign io_out_valid = ~io_hazard_in_stall; // @[2_Decode.scala 181:21]
  assign io_out_bits_isBranch = ctrlUnit_io_out_isBranch; // @[2_Decode.scala 150:29]
  assign io_out_bits_isJump = ctrlUnit_io_out_isJump; // @[2_Decode.scala 151:29]
  assign io_out_bits_resultSrc = ctrlUnit_io_out_resultSrc; // @[2_Decode.scala 152:29]
  assign io_out_bits_lsuOp = ctrlUnit_io_out_lsuOp; // @[2_Decode.scala 153:29]
  assign io_out_bits_aluOpSel = ctrlUnit_io_out_aluOpSel; // @[2_Decode.scala 154:29]
  assign io_out_bits_immSign = ctrlUnit_io_out_immSign; // @[2_Decode.scala 157:29]
  assign io_out_bits_regWrEn = ctrlUnit_io_out_regWrEn; // @[2_Decode.scala 156:29]
  assign io_out_bits_pcAddReg = ctrlUnit_io_out_pcAddReg; // @[2_Decode.scala 155:29]
  assign io_out_bits_pcNext4 = stageReg_pcNext4; // @[2_Decode.scala 173:29]
  assign io_out_bits_aluIn1 = 4'h8 == ctrlUnit_io_out_aluSrc1 ? 32'h4 : _io_out_bits_aluIn1_T_9; // @[Mux.scala 81:58]
  assign io_out_bits_aluIn2 = 4'h8 == ctrlUnit_io_out_aluSrc2 ? 32'h4 : _io_out_bits_aluIn2_T_9; // @[Mux.scala 81:58]
  assign io_out_bits_aluIn1IsReg = ctrlUnit_io_out_aluSrc1 == 4'h1 | ctrlUnit_io_out_aluSrc1 == 4'h2; // @[2_Decode.scala 168:54]
  assign io_out_bits_aluIn2IsReg = ctrlUnit_io_out_aluSrc2 == 4'h1 | ctrlUnit_io_out_aluSrc2 == 4'h2; // @[2_Decode.scala 169:54]
  assign io_out_bits_imm = immGen_io_imm; // @[2_Decode.scala 146:25 96:25]
  assign io_out_bits_data2 = io_regfile_rdata2; // @[2_Decode.scala 140:21 98:29]
  assign io_out_bits_excType = ctrlUnit_io_out_excType; // @[2_Decode.scala 162:29]
  assign io_out_bits_csrOp = ctrlUnit_io_out_csrOp; // @[2_Decode.scala 161:29]
  assign io_out_bits_instState_commit = io_ctrl_flush ? 1'h0 : stageReg_instState_commit; // @[2_Decode.scala 175:40]
  assign io_out_bits_instState_pc = stageReg_instState_pc; // @[2_Decode.scala 174:29]
  assign io_out_bits_instState_inst = stageReg_instState_inst; // @[2_Decode.scala 174:29]
  assign io_hazard_out_rs1 = stageReg_instState_inst[19:15]; // @[util.scala 72:31]
  assign io_hazard_out_rs2 = stageReg_instState_inst[24:20]; // @[util.scala 73:31]
  assign io_regfile_rs1 = stageReg_instState_inst[19:15]; // @[util.scala 72:31]
  assign io_regfile_rs2 = stageReg_instState_inst[24:20]; // @[util.scala 73:31]
  assign ctrlUnit_io_in_inst = stageReg_instState_inst; // @[2_Decode.scala 134:25]
  assign immGen_io_inst = stageReg_instState_inst; // @[2_Decode.scala 143:25]
  assign immGen_io_immSrc = ctrlUnit_io_out_immSrc; // @[2_Decode.scala 144:25]
  assign immGen_io_immSign = ctrlUnit_io_out_immSign; // @[2_Decode.scala 145:25]
  always @(posedge clock) begin
    if (reset) begin // @[2_Decode.scala 82:27]
      stageReg_pcNext4 <= 32'h0; // @[2_Decode.scala 82:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[2_Decode.scala 90:27]
      stageReg_pcNext4 <= 32'h0; // @[2_Decode.scala 90:38]
    end else if (decodeLatch) begin // @[2_Decode.scala 83:23]
      if (io_in_bits_instState_commit) begin // @[2_Decode.scala 84:24]
        stageReg_pcNext4 <= io_in_bits_pcNext4;
      end else begin
        stageReg_pcNext4 <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[2_Decode.scala 85:28]
      stageReg_pcNext4 <= 32'h0; // @[2_Decode.scala 86:18]
    end
    if (reset) begin // @[2_Decode.scala 82:27]
      stageReg_instState_commit <= 1'h0; // @[2_Decode.scala 82:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[2_Decode.scala 90:27]
      stageReg_instState_commit <= 1'h0; // @[2_Decode.scala 90:38]
    end else if (decodeLatch) begin // @[2_Decode.scala 83:23]
      stageReg_instState_commit <= io_in_bits_instState_commit; // @[2_Decode.scala 84:18]
    end else if (_io_in_ready_T_2) begin // @[2_Decode.scala 85:28]
      stageReg_instState_commit <= 1'h0; // @[2_Decode.scala 86:18]
    end
    if (reset) begin // @[2_Decode.scala 82:27]
      stageReg_instState_pc <= 32'h0; // @[2_Decode.scala 82:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[2_Decode.scala 90:27]
      stageReg_instState_pc <= 32'h0; // @[2_Decode.scala 90:38]
    end else if (decodeLatch) begin // @[2_Decode.scala 83:23]
      if (io_in_bits_instState_commit) begin // @[2_Decode.scala 84:24]
        stageReg_instState_pc <= io_in_bits_instState_pc;
      end else begin
        stageReg_instState_pc <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[2_Decode.scala 85:28]
      stageReg_instState_pc <= 32'h0; // @[2_Decode.scala 86:18]
    end
    if (reset) begin // @[2_Decode.scala 82:27]
      stageReg_instState_inst <= 32'h0; // @[2_Decode.scala 82:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[2_Decode.scala 90:27]
      stageReg_instState_inst <= 32'h0; // @[2_Decode.scala 90:38]
    end else if (decodeLatch) begin // @[2_Decode.scala 83:23]
      if (io_in_bits_instState_commit) begin // @[2_Decode.scala 84:24]
        stageReg_instState_inst <= io_in_bits_instState_inst;
      end else begin
        stageReg_instState_inst <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[2_Decode.scala 85:28]
      stageReg_instState_inst <= 32'h0; // @[2_Decode.scala 86:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stageReg_pcNext4 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stageReg_instState_commit = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  stageReg_instState_pc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  stageReg_instState_inst = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  input  [3:0]  io_opSel,
  output [31:0] io_out,
  output        io_zero
);
  wire [31:0] _sum_T_2 = 32'h0 - io_in2; // @[Alu.scala 25:41]
  wire [31:0] _sum_T_3 = io_opSel[0] ? _sum_T_2 : io_in2; // @[Alu.scala 25:27]
  wire [31:0] sum = io_in1 + _sum_T_3; // @[Alu.scala 25:22]
  wire [4:0] shamt = io_in2[4:0]; // @[Alu.scala 28:23]
  wire [31:0] _shiftr_T_1 = io_in1 >> shamt; // @[Alu.scala 30:32]
  wire [31:0] _shiftr_T_4 = $signed(io_in1) >>> shamt; // @[Alu.scala 31:49]
  wire [31:0] shiftr = io_opSel[1] ? _shiftr_T_1 : _shiftr_T_4; // @[Alu.scala 29:21]
  wire [62:0] _GEN_5 = {{31'd0}, io_in1}; // @[Alu.scala 33:25]
  wire [62:0] shiftl = _GEN_5 << shamt; // @[Alu.scala 33:25]
  wire [31:0] _shout_T_3 = io_opSel == 4'hb | io_opSel == 4'hc ? shiftr : 32'h0; // @[Alu.scala 34:20]
  wire [62:0] _shout_T_5 = io_opSel == 4'ha ? shiftl : 63'h0; // @[Alu.scala 35:20]
  wire [62:0] _GEN_2 = {{31'd0}, _shout_T_3}; // @[Alu.scala 34:80]
  wire [62:0] shout = _GEN_2 | _shout_T_5; // @[Alu.scala 34:80]
  wire [31:0] _logic_T = io_in1 & io_in2; // @[Alu.scala 40:40]
  wire [31:0] _logic_T_1 = io_in1 | io_in2; // @[Alu.scala 41:40]
  wire [31:0] _logic_T_2 = io_in1 ^ io_in2; // @[Alu.scala 42:40]
  wire [31:0] _logic_T_4 = 4'h2 == io_opSel ? _logic_T : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _logic_T_6 = 4'h3 == io_opSel ? _logic_T_1 : _logic_T_4; // @[Mux.scala 81:58]
  wire [31:0] logic_ = 4'h4 == io_opSel ? _logic_T_2 : _logic_T_6; // @[Mux.scala 81:58]
  wire  _cmp_T_2 = $signed(io_in1) < $signed(io_in2); // @[Alu.scala 48:48]
  wire  _cmp_T_3 = io_in1 < io_in2; // @[Alu.scala 49:41]
  wire  _cmp_T_4 = io_in1 == io_in2; // @[Alu.scala 50:41]
  wire  _cmp_T_5 = io_in1 != io_in2; // @[Alu.scala 51:41]
  wire  _cmp_T_8 = $signed(io_in1) >= $signed(io_in2); // @[Alu.scala 52:48]
  wire  _cmp_T_9 = io_in1 >= io_in2; // @[Alu.scala 53:42]
  wire  _cmp_T_13 = 4'h9 == io_opSel ? _cmp_T_3 : 4'h8 == io_opSel & _cmp_T_2; // @[Mux.scala 81:58]
  wire  _cmp_T_15 = 4'h5 == io_opSel ? _cmp_T_4 : _cmp_T_13; // @[Mux.scala 81:58]
  wire  _cmp_T_17 = 4'h6 == io_opSel ? _cmp_T_5 : _cmp_T_15; // @[Mux.scala 81:58]
  wire  _cmp_T_19 = 4'h7 == io_opSel ? _cmp_T_8 : _cmp_T_17; // @[Mux.scala 81:58]
  wire  cmp = 4'hf == io_opSel ? _cmp_T_9 : _cmp_T_19; // @[Mux.scala 81:58]
  wire [31:0] _GEN_3 = {{31'd0}, cmp}; // @[Alu.scala 62:66]
  wire [31:0] _io_out_T_3 = _GEN_3 | logic_; // @[Alu.scala 62:66]
  wire [62:0] _GEN_4 = {{31'd0}, _io_out_T_3}; // @[Alu.scala 62:74]
  wire [62:0] _io_out_T_4 = _GEN_4 | shout; // @[Alu.scala 62:74]
  wire [62:0] _io_out_T_5 = io_opSel == 4'h0 | io_opSel == 4'h1 ? {{31'd0}, sum} : _io_out_T_4; // @[Alu.scala 62:22]
  wire [62:0] _GEN_0 = io_opSel == 4'he ? {{31'd0}, io_in2} : _io_out_T_5; // @[Alu.scala 59:33 60:16 62:16]
  wire [62:0] _GEN_1 = io_opSel == 4'hd ? {{31'd0}, io_in1} : _GEN_0; // @[Alu.scala 57:27 58:16]
  assign io_out = _GEN_1[31:0];
  assign io_zero = 4'hf == io_opSel ? _cmp_T_9 : _cmp_T_19; // @[Mux.scala 81:58]
endmodule
module Execute(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_isBranch,
  input         io_in_bits_isJump,
  input  [1:0]  io_in_bits_resultSrc,
  input  [4:0]  io_in_bits_lsuOp,
  input  [3:0]  io_in_bits_aluOpSel,
  input         io_in_bits_immSign,
  input         io_in_bits_regWrEn,
  input         io_in_bits_pcAddReg,
  input  [31:0] io_in_bits_pcNext4,
  input  [31:0] io_in_bits_aluIn1,
  input  [31:0] io_in_bits_aluIn2,
  input         io_in_bits_aluIn1IsReg,
  input         io_in_bits_aluIn2IsReg,
  input  [31:0] io_in_bits_imm,
  input  [31:0] io_in_bits_data2,
  input  [3:0]  io_in_bits_excType,
  input  [2:0]  io_in_bits_csrOp,
  input         io_in_bits_instState_commit,
  input  [31:0] io_in_bits_instState_pc,
  input  [31:0] io_in_bits_instState_inst,
  input         io_out_memory_ready,
  output        io_out_memory_valid,
  output [1:0]  io_out_memory_bits_resultSrc,
  output [4:0]  io_out_memory_bits_lsuOp,
  output        io_out_memory_bits_regWrEn,
  output [31:0] io_out_memory_bits_aluOut,
  output [31:0] io_out_memory_bits_data2,
  output [31:0] io_out_memory_bits_pcNext4,
  output [2:0]  io_out_memory_bits_csrOp,
  output        io_out_memory_bits_csrWrEn,
  output        io_out_memory_bits_csrValid,
  output [31:0] io_out_memory_bits_csrRdData,
  output [31:0] io_out_memory_bits_csrWrData,
  output [31:0] io_out_memory_bits_csrAddr,
  output [3:0]  io_out_memory_bits_excType,
  output        io_out_memory_bits_instState_commit,
  output [31:0] io_out_memory_bits_instState_pc,
  output [31:0] io_out_memory_bits_instState_inst,
  output        io_out_fetch_bits_brTaken,
  output [31:0] io_out_fetch_bits_targetAddr,
  output [4:0]  io_hazard_out_rs1,
  output [4:0]  io_hazard_out_rs2,
  output [1:0]  io_hazard_out_resultSrc,
  output [4:0]  io_hazard_out_rd,
  input  [1:0]  io_hazard_in_aluSrc1,
  input  [1:0]  io_hazard_in_aluSrc2,
  input  [31:0] io_hazard_in_rdValM,
  input  [31:0] io_hazard_in_rdValW,
  input         io_ctrl_flush,
  output [2:0]  io_csrRead_op,
  input         io_csrRead_valid,
  output [11:0] io_csrRead_addr,
  input  [31:0] io_csrRead_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] alu_io_in1; // @[3_Execute.scala 102:29]
  wire [31:0] alu_io_in2; // @[3_Execute.scala 102:29]
  wire [3:0] alu_io_opSel; // @[3_Execute.scala 102:29]
  wire [31:0] alu_io_out; // @[3_Execute.scala 102:29]
  wire  alu_io_zero; // @[3_Execute.scala 102:29]
  wire  _io_in_ready_T_2 = io_out_memory_ready & io_out_memory_valid; // @[Decoupled.scala 51:35]
  wire  executeLatch = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  reg  stageReg_isBranch; // @[3_Execute.scala 89:27]
  reg  stageReg_isJump; // @[3_Execute.scala 89:27]
  reg [1:0] stageReg_resultSrc; // @[3_Execute.scala 89:27]
  reg [4:0] stageReg_lsuOp; // @[3_Execute.scala 89:27]
  reg [3:0] stageReg_aluOpSel; // @[3_Execute.scala 89:27]
  reg  stageReg_immSign; // @[3_Execute.scala 89:27]
  reg  stageReg_regWrEn; // @[3_Execute.scala 89:27]
  reg  stageReg_pcAddReg; // @[3_Execute.scala 89:27]
  reg [31:0] stageReg_pcNext4; // @[3_Execute.scala 89:27]
  reg [31:0] stageReg_aluIn1; // @[3_Execute.scala 89:27]
  reg [31:0] stageReg_aluIn2; // @[3_Execute.scala 89:27]
  reg  stageReg_aluIn1IsReg; // @[3_Execute.scala 89:27]
  reg  stageReg_aluIn2IsReg; // @[3_Execute.scala 89:27]
  reg [31:0] stageReg_imm; // @[3_Execute.scala 89:27]
  reg [31:0] stageReg_data2; // @[3_Execute.scala 89:27]
  reg [3:0] stageReg_excType; // @[3_Execute.scala 89:27]
  reg [2:0] stageReg_csrOp; // @[3_Execute.scala 89:27]
  reg  stageReg_instState_commit; // @[3_Execute.scala 89:27]
  reg [31:0] stageReg_instState_pc; // @[3_Execute.scala 89:27]
  reg [31:0] stageReg_instState_inst; // @[3_Execute.scala 89:27]
  wire [31:0] _hazardData1_T_3 = 2'h1 == io_hazard_in_aluSrc1 ? io_hazard_in_rdValM : stageReg_aluIn1; // @[Mux.scala 81:58]
  wire [31:0] hazardData1 = 2'h2 == io_hazard_in_aluSrc1 ? io_hazard_in_rdValW : _hazardData1_T_3; // @[Mux.scala 81:58]
  wire [31:0] _hazardData2_T_3 = 2'h1 == io_hazard_in_aluSrc2 ? io_hazard_in_rdValM : stageReg_aluIn2; // @[Mux.scala 81:58]
  wire [31:0] hazardData2 = 2'h2 == io_hazard_in_aluSrc2 ? io_hazard_in_rdValW : _hazardData2_T_3; // @[Mux.scala 81:58]
  wire  aluZero = alu_io_zero; // @[3_Execute.scala 134:18 98:23]
  wire [31:0] _io_out_fetch_bits_targetAddr_T_5 = $signed(stageReg_imm) + $signed(stageReg_instState_pc); // @[3_Execute.scala 140:102]
  wire [31:0] _io_out_fetch_bits_targetAddr_T_7 = stageReg_imm + stageReg_instState_pc; // @[3_Execute.scala 141:62]
  wire [31:0] _io_out_fetch_bits_targetAddr_T_8 = stageReg_immSign ? _io_out_fetch_bits_targetAddr_T_5 :
    _io_out_fetch_bits_targetAddr_T_7; // @[3_Execute.scala 139:48]
  wire [31:0] _io_out_memory_bits_data2_T_3 = io_hazard_in_aluSrc2 == 2'h2 ? io_hazard_in_rdValW : stageReg_data2; // @[3_Execute.scala 155:52]
  wire [31:0] _io_out_memory_bits_data2_T_4 = io_hazard_in_aluSrc2 == 2'h1 ? io_hazard_in_rdValM :
    _io_out_memory_bits_data2_T_3; // @[3_Execute.scala 153:48]
  wire [11:0] csrAddr = stageReg_instState_inst[31:20]; // @[util.scala 78:36]
  ALU alu ( // @[3_Execute.scala 102:29]
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_opSel(alu_io_opSel),
    .io_out(alu_io_out),
    .io_zero(alu_io_zero)
  );
  assign io_in_ready = io_in_valid & _io_in_ready_T_2; // @[3_Execute.scala 87:43]
  assign io_out_memory_valid = 1'h1; // @[3_Execute.scala 190:39]
  assign io_out_memory_bits_resultSrc = stageReg_resultSrc; // @[3_Execute.scala 148:37]
  assign io_out_memory_bits_lsuOp = stageReg_lsuOp; // @[3_Execute.scala 149:37]
  assign io_out_memory_bits_regWrEn = stageReg_regWrEn; // @[3_Execute.scala 150:37]
  assign io_out_memory_bits_aluOut = alu_io_out; // @[3_Execute.scala 147:37]
  assign io_out_memory_bits_data2 = io_hazard_in_aluSrc2 == 2'h0 ? stageReg_data2 : _io_out_memory_bits_data2_T_4; // @[3_Execute.scala 151:43]
  assign io_out_memory_bits_pcNext4 = stageReg_pcNext4; // @[3_Execute.scala 161:37]
  assign io_out_memory_bits_csrOp = stageReg_csrOp; // @[3_Execute.scala 168:35]
  assign io_out_memory_bits_csrWrEn = stageReg_csrOp != 3'h0 & io_csrRead_valid; // @[3_Execute.scala 169:65]
  assign io_out_memory_bits_csrValid = io_csrRead_valid; // @[3_Execute.scala 170:35]
  assign io_out_memory_bits_csrRdData = io_csrRead_data; // @[3_Execute.scala 171:35]
  assign io_out_memory_bits_csrWrData = stageReg_aluIn1IsReg ? hazardData1 : stageReg_aluIn1; // @[3_Execute.scala 118:27]
  assign io_out_memory_bits_csrAddr = {{20'd0}, csrAddr}; // @[3_Execute.scala 173:35]
  assign io_out_memory_bits_excType = stageReg_excType; // @[3_Execute.scala 174:35]
  assign io_out_memory_bits_instState_commit = io_ctrl_flush ? 1'h0 : stageReg_instState_commit; // @[3_Execute.scala 187:47]
  assign io_out_memory_bits_instState_pc = stageReg_instState_pc; // @[3_Execute.scala 186:35]
  assign io_out_memory_bits_instState_inst = stageReg_instState_inst; // @[3_Execute.scala 186:35]
  assign io_out_fetch_bits_brTaken = (stageReg_isBranch & aluZero | stageReg_isJump) & stageReg_instState_commit; // @[3_Execute.scala 137:94]
  assign io_out_fetch_bits_targetAddr = stageReg_pcAddReg ? alu_io_out : _io_out_fetch_bits_targetAddr_T_8; // @[3_Execute.scala 138:43]
  assign io_hazard_out_rs1 = stageReg_instState_inst[19:15]; // @[util.scala 72:31]
  assign io_hazard_out_rs2 = stageReg_instState_inst[24:20]; // @[util.scala 73:31]
  assign io_hazard_out_resultSrc = stageReg_resultSrc; // @[3_Execute.scala 182:35]
  assign io_hazard_out_rd = stageReg_instState_inst[11:7]; // @[util.scala 71:31]
  assign io_csrRead_op = stageReg_csrOp; // @[3_Execute.scala 167:35]
  assign io_csrRead_addr = stageReg_instState_inst[31:20]; // @[util.scala 78:36]
  assign alu_io_in1 = stageReg_aluIn1IsReg ? hazardData1 : stageReg_aluIn1; // @[3_Execute.scala 118:27]
  assign alu_io_in2 = stageReg_aluIn2IsReg ? hazardData2 : stageReg_aluIn2; // @[3_Execute.scala 120:27]
  assign alu_io_opSel = stageReg_aluOpSel; // @[3_Execute.scala 133:18]
  always @(posedge clock) begin
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_isBranch <= 1'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_isBranch <= 1'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      stageReg_isBranch <= io_in_bits_instState_commit & io_in_bits_isBranch; // @[3_Execute.scala 91:18]
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_isBranch <= 1'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_isJump <= 1'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_isJump <= 1'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      stageReg_isJump <= io_in_bits_instState_commit & io_in_bits_isJump; // @[3_Execute.scala 91:18]
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_isJump <= 1'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_resultSrc <= 2'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_resultSrc <= 2'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_resultSrc <= io_in_bits_resultSrc;
      end else begin
        stageReg_resultSrc <= 2'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_resultSrc <= 2'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_lsuOp <= 5'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_lsuOp <= 5'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_lsuOp <= io_in_bits_lsuOp;
      end else begin
        stageReg_lsuOp <= 5'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_lsuOp <= 5'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_aluOpSel <= 4'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_aluOpSel <= 4'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_aluOpSel <= io_in_bits_aluOpSel;
      end else begin
        stageReg_aluOpSel <= 4'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_aluOpSel <= 4'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_immSign <= 1'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_immSign <= 1'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      stageReg_immSign <= io_in_bits_instState_commit & io_in_bits_immSign; // @[3_Execute.scala 91:18]
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_immSign <= 1'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_regWrEn <= 1'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_regWrEn <= 1'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      stageReg_regWrEn <= io_in_bits_instState_commit & io_in_bits_regWrEn; // @[3_Execute.scala 91:18]
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_regWrEn <= 1'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_pcAddReg <= 1'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_pcAddReg <= 1'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      stageReg_pcAddReg <= io_in_bits_instState_commit & io_in_bits_pcAddReg; // @[3_Execute.scala 91:18]
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_pcAddReg <= 1'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_pcNext4 <= 32'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_pcNext4 <= 32'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_pcNext4 <= io_in_bits_pcNext4;
      end else begin
        stageReg_pcNext4 <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_pcNext4 <= 32'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_aluIn1 <= 32'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_aluIn1 <= 32'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_aluIn1 <= io_in_bits_aluIn1;
      end else begin
        stageReg_aluIn1 <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_aluIn1 <= 32'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_aluIn2 <= 32'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_aluIn2 <= 32'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_aluIn2 <= io_in_bits_aluIn2;
      end else begin
        stageReg_aluIn2 <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_aluIn2 <= 32'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_aluIn1IsReg <= 1'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_aluIn1IsReg <= 1'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      stageReg_aluIn1IsReg <= io_in_bits_instState_commit & io_in_bits_aluIn1IsReg; // @[3_Execute.scala 91:18]
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_aluIn1IsReg <= 1'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_aluIn2IsReg <= 1'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_aluIn2IsReg <= 1'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      stageReg_aluIn2IsReg <= io_in_bits_instState_commit & io_in_bits_aluIn2IsReg; // @[3_Execute.scala 91:18]
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_aluIn2IsReg <= 1'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_imm <= 32'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_imm <= 32'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_imm <= io_in_bits_imm;
      end else begin
        stageReg_imm <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_imm <= 32'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_data2 <= 32'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_data2 <= 32'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_data2 <= io_in_bits_data2;
      end else begin
        stageReg_data2 <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_data2 <= 32'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_excType <= 4'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_excType <= 4'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_excType <= io_in_bits_excType;
      end else begin
        stageReg_excType <= 4'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_excType <= 4'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_csrOp <= 3'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_csrOp <= 3'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_csrOp <= io_in_bits_csrOp;
      end else begin
        stageReg_csrOp <= 3'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_csrOp <= 3'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_instState_commit <= 1'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_instState_commit <= 1'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      stageReg_instState_commit <= io_in_bits_instState_commit; // @[3_Execute.scala 91:18]
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_instState_commit <= 1'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_instState_pc <= 32'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_instState_pc <= 32'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_instState_pc <= io_in_bits_instState_pc;
      end else begin
        stageReg_instState_pc <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_instState_pc <= 32'h0; // @[3_Execute.scala 93:18]
    end
    if (reset) begin // @[3_Execute.scala 89:27]
      stageReg_instState_inst <= 32'h0; // @[3_Execute.scala 89:27]
    end else if (io_ctrl_flush) begin // @[3_Execute.scala 96:27]
      stageReg_instState_inst <= 32'h0; // @[3_Execute.scala 96:38]
    end else if (executeLatch) begin // @[3_Execute.scala 90:24]
      if (io_in_bits_instState_commit) begin // @[3_Execute.scala 91:24]
        stageReg_instState_inst <= io_in_bits_instState_inst;
      end else begin
        stageReg_instState_inst <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[3_Execute.scala 92:35]
      stageReg_instState_inst <= 32'h0; // @[3_Execute.scala 93:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stageReg_isBranch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stageReg_isJump = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  stageReg_resultSrc = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  stageReg_lsuOp = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  stageReg_aluOpSel = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  stageReg_immSign = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  stageReg_regWrEn = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  stageReg_pcAddReg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  stageReg_pcNext4 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  stageReg_aluIn1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  stageReg_aluIn2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  stageReg_aluIn1IsReg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  stageReg_aluIn2IsReg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  stageReg_imm = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  stageReg_data2 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  stageReg_excType = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  stageReg_csrOp = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  stageReg_instState_commit = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  stageReg_instState_pc = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  stageReg_instState_inst = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSU_1(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [31:0] io_req_bits_addr,
  input  [31:0] io_req_bits_wdata,
  input  [4:0]  io_req_bits_lsuOp,
  output        io_resp_valid,
  output [31:0] io_resp_bits_rdata,
  input         io_cache_read_req_ready,
  output        io_cache_read_req_valid,
  output [31:0] io_cache_read_req_bits_addr,
  output        io_cache_read_resp_ready,
  input         io_cache_read_resp_valid,
  input  [31:0] io_cache_read_resp_bits_data,
  input         io_cache_write_req_ready,
  output        io_cache_write_req_valid,
  output [31:0] io_cache_write_req_bits_addr,
  output [31:0] io_cache_write_req_bits_data,
  output [3:0]  io_cache_write_req_bits_mask,
  output        io_cache_write_resp_ready,
  input         io_cache_write_resp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg  s0_full; // @[LSU.scala 206:26]
  wire  s0_latch = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  wire  _s0_valid_T = io_cache_read_req_ready & io_cache_read_req_valid; // @[Decoupled.scala 51:35]
  reg  s0_valid_holdReg; // @[Reg.scala 19:16]
  wire  _s0_valid_T_1 = _s0_valid_T | s0_valid_holdReg; // @[util.scala 26:12]
  reg [4:0] s0_reqReg_lsuOp; // @[Reg.scala 19:16]
  wire [4:0] s0_req_lsuOp = s0_latch ? io_req_bits_lsuOp : s0_reqReg_lsuOp; // @[LSU.scala 211:21]
  wire  _T_7 = 5'h1 == s0_req_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_9 = 5'h2 == s0_req_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_11 = 5'h3 == s0_req_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_13 = 5'h4 == s0_req_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_15 = 5'h5 == s0_req_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_17 = 5'h6 == s0_req_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_19 = 5'h7 == s0_req_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_21 = 5'h8 == s0_req_lsuOp; // @[Lookup.scala 31:38]
  wire  load = _T_7 | (_T_9 | (_T_11 | (_T_13 | _T_15))); // @[Lookup.scala 34:39]
  wire  _s0_valid_T_3 = io_cache_write_req_ready & io_cache_write_req_valid; // @[Decoupled.scala 51:35]
  reg  s0_valid_holdReg_1; // @[Reg.scala 19:16]
  wire  _s0_valid_T_4 = _s0_valid_T_3 | s0_valid_holdReg_1; // @[util.scala 26:12]
  wire  _T_36 = _T_15 ? 1'h0 : _T_17 | (_T_19 | _T_21); // @[Lookup.scala 34:39]
  wire  _T_37 = _T_13 ? 1'h0 : _T_36; // @[Lookup.scala 34:39]
  wire  _T_38 = _T_11 ? 1'h0 : _T_37; // @[Lookup.scala 34:39]
  wire  _T_39 = _T_9 ? 1'h0 : _T_38; // @[Lookup.scala 34:39]
  wire  wen = _T_7 ? 1'h0 : _T_39; // @[Lookup.scala 34:39]
  wire  s0_valid = _s0_valid_T_1 & load | _s0_valid_T_4 & wen; // @[LSU.scala 265:73]
  reg  s1_full; // @[LSU.scala 272:26]
  wire  s1_ready = ~s1_full; // @[LSU.scala 279:17]
  wire  s0_fire = s0_valid & s1_ready; // @[LSU.scala 208:28]
  reg [31:0] s0_reqReg_addr; // @[Reg.scala 19:16]
  reg [31:0] s0_reqReg_wdata; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = s0_latch ? io_req_bits_addr : s0_reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_1 = s0_latch ? io_req_bits_wdata : s0_reqReg_wdata; // @[Reg.scala 19:16 20:{18,22}]
  wire [1:0] s0_offset = _GEN_0[1:0]; // @[LSU.scala 212:32]
  wire  _GEN_4 = s0_full & s0_fire ? 1'h0 : s0_full; // @[LSU.scala 206:26 217:{35,45}]
  wire  _GEN_5 = s0_latch & ~(s0_req_lsuOp == 5'h0 | s0_req_lsuOp == 5'h14) | _GEN_4; // @[LSU.scala 216:{80,90}]
  wire  en = _T_7 | (_T_9 | (_T_11 | (_T_13 | (_T_15 | (_T_17 | (_T_19 | _T_21)))))); // @[Lookup.scala 34:39]
  wire [1:0] _T_49 = _T_21 ? 2'h2 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _T_50 = _T_19 ? 2'h1 : _T_49; // @[Lookup.scala 34:39]
  wire [1:0] _T_51 = _T_17 ? 2'h0 : _T_50; // @[Lookup.scala 34:39]
  wire [1:0] _T_52 = _T_15 ? 2'h1 : _T_51; // @[Lookup.scala 34:39]
  wire [1:0] _T_53 = _T_13 ? 2'h0 : _T_52; // @[Lookup.scala 34:39]
  wire [1:0] _T_54 = _T_11 ? 2'h2 : _T_53; // @[Lookup.scala 34:39]
  wire [1:0] _T_55 = _T_9 ? 2'h1 : _T_54; // @[Lookup.scala 34:39]
  wire [1:0] width = _T_7 ? 2'h0 : _T_55; // @[Lookup.scala 34:39]
  wire  signed_ = _T_7 | (_T_9 | (_T_11 | _T_37)); // @[Lookup.scala 34:39]
  wire  _s0_reqSend_T_2 = _s0_valid_T | _s0_valid_T_3; // @[LSU.scala 243:72]
  reg  s0_reqSend; // @[Reg.scala 35:20]
  wire  _GEN_8 = _s0_reqSend_T_2 | s0_reqSend; // @[Reg.scala 36:18 35:20 36:22]
  wire  _io_cache_read_req_valid_T_1 = ~s0_reqSend; // @[LSU.scala 245:51]
  wire [4:0] _io_cache_write_req_bits_data_T = {s0_offset, 3'h0}; // @[LSU.scala 250:64]
  wire [62:0] _GEN_2 = {{31'd0}, _GEN_1}; // @[LSU.scala 250:50]
  wire [62:0] _io_cache_write_req_bits_data_T_1 = _GEN_2 << _io_cache_write_req_bits_data_T; // @[LSU.scala 250:50]
  wire [3:0] _s0_storeMask_T_1 = 4'h1 << s0_offset; // @[OneHot.scala 57:35]
  wire [2:0] _s0_storeMask_T_6 = 2'h1 == s0_offset ? 3'h6 : 3'h3; // @[Mux.scala 81:58]
  wire [3:0] _s0_storeMask_T_8 = 2'h2 == s0_offset ? 4'hc : {{1'd0}, _s0_storeMask_T_6}; // @[Mux.scala 81:58]
  wire [3:0] _s0_storeMask_T_10 = 2'h0 == width ? _s0_storeMask_T_1 : 4'hf; // @[Mux.scala 81:58]
  wire [3:0] _s0_storeMask_T_12 = 2'h1 == width ? _s0_storeMask_T_8 : _s0_storeMask_T_10; // @[Mux.scala 81:58]
  reg  s1_signed; // @[Reg.scala 19:16]
  reg [1:0] s1_width; // @[Reg.scala 19:16]
  reg [1:0] s1_offset; // @[Reg.scala 19:16]
  wire  _s1_loadRespValid_T = io_cache_read_resp_ready & io_cache_read_resp_valid; // @[Decoupled.scala 51:35]
  reg  s1_loadRespValid_holdReg; // @[Reg.scala 19:16]
  wire  s1_loadRespValid = _s1_loadRespValid_T ? io_cache_read_resp_valid : s1_loadRespValid_holdReg; // @[util.scala 26:12]
  wire  _s1_storeRespValid_T = io_cache_write_resp_ready & io_cache_write_resp_valid; // @[Decoupled.scala 51:35]
  reg  s1_storeRespValid_holdReg; // @[Reg.scala 19:16]
  wire  s1_storeRespValid = _s1_storeRespValid_T ? io_cache_write_resp_valid : s1_storeRespValid_holdReg; // @[util.scala 26:12]
  wire  s1_fire = s1_full & (s1_loadRespValid | s1_storeRespValid); // @[LSU.scala 306:25]
  wire  _GEN_17 = s1_full & s1_fire ? 1'h0 : s1_full; // @[LSU.scala 272:26 281:{35,45}]
  wire  _GEN_18 = s0_fire | _GEN_17; // @[LSU.scala 280:{20,30}]
  reg [31:0] s1_loadResp_holdReg_data; // @[Reg.scala 19:16]
  wire [31:0] _GEN_21 = _s1_loadRespValid_T ? io_cache_read_resp_bits_data : s1_loadResp_holdReg_data; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _s1_loadData_T_2 = {8'h0,_GEN_21[31:8]}; // @[Cat.scala 33:92]
  wire [31:0] _s1_loadData_T_5 = {16'h0,_GEN_21[31:16]}; // @[Cat.scala 33:92]
  wire [31:0] _s1_loadData_T_8 = {24'h0,_GEN_21[31:24]}; // @[Cat.scala 33:92]
  wire [31:0] _s1_loadData_T_10 = 2'h1 == s1_offset ? _s1_loadData_T_2 : _GEN_21; // @[Mux.scala 81:58]
  wire [31:0] _s1_loadData_T_12 = 2'h2 == s1_offset ? _s1_loadData_T_5 : _s1_loadData_T_10; // @[Mux.scala 81:58]
  wire [31:0] s1_loadData = 2'h3 == s1_offset ? _s1_loadData_T_8 : _s1_loadData_T_12; // @[Mux.scala 81:58]
  wire [7:0] _io_resp_bits_rdata_T_1 = s1_loadData[7:0]; // @[LSU.scala 300:85]
  wire  io_resp_bits_rdata_signBit = _io_resp_bits_rdata_T_1[7]; // @[util.scala 42:27]
  wire [5:0] io_resp_bits_rdata_out_lo_lo = {io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,
    io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit}; // @[Cat.scala 33:92]
  wire [11:0] io_resp_bits_rdata_out_lo = {io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,
    io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,
    io_resp_bits_rdata_out_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] _io_resp_bits_rdata_out_T_1 = s1_loadData[7:0]; // @[util.scala 46:75]
  wire [31:0] io_resp_bits_rdata_out = {io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit
    ,io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,io_resp_bits_rdata_signBit,io_resp_bits_rdata_out_lo_lo,
    io_resp_bits_rdata_out_lo,_io_resp_bits_rdata_out_T_1}; // @[Cat.scala 33:92]
  wire [31:0] io_resp_bits_rdata_out_1 = {{24'd0}, s1_loadData[7:0]}; // @[util.scala 62:36]
  wire [31:0] _io_resp_bits_rdata_T_3 = s1_signed ? io_resp_bits_rdata_out : io_resp_bits_rdata_out_1; // @[LSU.scala 300:48]
  wire [15:0] _io_resp_bits_rdata_T_5 = s1_loadData[15:0]; // @[LSU.scala 301:86]
  wire  io_resp_bits_rdata_signBit_1 = _io_resp_bits_rdata_T_5[15]; // @[util.scala 42:27]
  wire [7:0] io_resp_bits_rdata_out_lo_1 = {io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1,
    io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1,
    io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1}; // @[Cat.scala 33:92]
  wire [15:0] _io_resp_bits_rdata_out_T_3 = s1_loadData[15:0]; // @[util.scala 46:75]
  wire [31:0] io_resp_bits_rdata_out_2 = {io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1,
    io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1,
    io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_signBit_1,io_resp_bits_rdata_out_lo_1,_io_resp_bits_rdata_out_T_3}; // @[Cat.scala 33:92]
  wire [31:0] io_resp_bits_rdata_out_3 = {{16'd0}, s1_loadData[15:0]}; // @[util.scala 62:36]
  wire [31:0] _io_resp_bits_rdata_T_7 = s1_signed ? io_resp_bits_rdata_out_2 : io_resp_bits_rdata_out_3; // @[LSU.scala 301:48]
  wire [31:0] _io_resp_bits_rdata_T_10 = 2'h3 == s1_offset ? _s1_loadData_T_8 : _s1_loadData_T_12; // @[util.scala 44:18]
  wire [31:0] _io_resp_bits_rdata_T_12 = s1_signed ? _io_resp_bits_rdata_T_10 : s1_loadData; // @[LSU.scala 302:48]
  wire [31:0] _io_resp_bits_rdata_T_14 = 2'h0 == s1_width ? _io_resp_bits_rdata_T_3 : s1_loadData; // @[Mux.scala 81:58]
  wire [31:0] _io_resp_bits_rdata_T_16 = 2'h1 == s1_width ? _io_resp_bits_rdata_T_7 : _io_resp_bits_rdata_T_14; // @[Mux.scala 81:58]
  wire  s0_en = en; // @[Lookup.scala 34:39]
  assign io_req_ready = ~s0_full; // @[LSU.scala 214:21]
  assign io_resp_valid = s1_full & (s1_loadRespValid | s1_storeRespValid); // @[LSU.scala 306:25]
  assign io_resp_bits_rdata = 2'h2 == s1_width ? _io_resp_bits_rdata_T_12 : _io_resp_bits_rdata_T_16; // @[Mux.scala 81:58]
  assign io_cache_read_req_valid = load & s0_full & ~s0_reqSend; // @[LSU.scala 245:48]
  assign io_cache_read_req_bits_addr = {_GEN_0[31:2],2'h0}; // @[Cat.scala 33:92]
  assign io_cache_read_resp_ready = 1'h1; // @[LSU.scala 283:30]
  assign io_cache_write_req_valid = wen & s0_full & _io_cache_read_req_valid_T_1; // @[LSU.scala 248:48]
  assign io_cache_write_req_bits_addr = {_GEN_0[31:2],2'h0}; // @[Cat.scala 33:92]
  assign io_cache_write_req_bits_data = _io_cache_write_req_bits_data_T_1[31:0]; // @[LSU.scala 250:34]
  assign io_cache_write_req_bits_mask = 2'h2 == width ? 4'hf : _s0_storeMask_T_12; // @[Mux.scala 81:58]
  assign io_cache_write_resp_ready = 1'h1; // @[LSU.scala 284:31]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 206:26]
      s0_full <= 1'h0; // @[LSU.scala 206:26]
    end else begin
      s0_full <= _GEN_5;
    end
    if (s0_fire) begin // @[util.scala 25:21]
      s0_valid_holdReg <= 1'h0; // @[util.scala 25:31]
    end else begin
      s0_valid_holdReg <= _s0_valid_T_1;
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_lsuOp <= io_req_bits_lsuOp; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[util.scala 25:21]
      s0_valid_holdReg_1 <= 1'h0; // @[util.scala 25:31]
    end else begin
      s0_valid_holdReg_1 <= _s0_valid_T_4;
    end
    if (reset) begin // @[LSU.scala 272:26]
      s1_full <= 1'h0; // @[LSU.scala 272:26]
    end else begin
      s1_full <= _GEN_18;
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_addr <= io_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_wdata <= io_req_bits_wdata; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      s0_reqSend <= 1'h0; // @[Reg.scala 35:20]
    end else if (s0_fire) begin // @[LSU.scala 244:19]
      s0_reqSend <= 1'h0; // @[LSU.scala 244:32]
    end else begin
      s0_reqSend <= _GEN_8;
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_signed <= signed_; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      if (_T_7) begin // @[Lookup.scala 34:39]
        s1_width <= 2'h0;
      end else if (_T_9) begin // @[Lookup.scala 34:39]
        s1_width <= 2'h1;
      end else if (_T_11) begin // @[Lookup.scala 34:39]
        s1_width <= 2'h2;
      end else begin
        s1_width <= _T_53;
      end
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_offset <= s0_offset; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[util.scala 25:21]
      s1_loadRespValid_holdReg <= 1'h0; // @[util.scala 25:31]
    end else if (_s1_loadRespValid_T) begin // @[util.scala 26:12]
      s1_loadRespValid_holdReg <= io_cache_read_resp_valid;
    end
    if (s0_fire) begin // @[util.scala 25:21]
      s1_storeRespValid_holdReg <= 1'h0; // @[util.scala 25:31]
    end else if (_s1_storeRespValid_T) begin // @[util.scala 26:12]
      s1_storeRespValid_holdReg <= io_cache_write_resp_valid;
    end
    if (s0_fire) begin // @[util.scala 25:21]
      s1_loadResp_holdReg_data <= 32'h0; // @[util.scala 25:31]
    end else if (_s1_loadRespValid_T) begin // @[Reg.scala 20:18]
      s1_loadResp_holdReg_data <= io_cache_read_resp_bits_data; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s0_valid_holdReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s0_reqReg_lsuOp = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  s0_valid_holdReg_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s1_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s0_reqReg_addr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  s0_reqReg_wdata = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  s0_reqSend = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s1_signed = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  s1_width = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  s1_offset = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  s1_loadRespValid_holdReg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  s1_storeRespValid_holdReg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  s1_loadResp_holdReg_data = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LoadPipe(
  input         clock,
  input         reset,
  output        io_load_req_ready,
  input         io_load_req_valid,
  input  [31:0] io_load_req_bits_addr,
  output        io_load_resp_valid,
  output [31:0] io_load_resp_bits_data,
  input         io_dir_req_ready,
  output        io_dir_req_valid,
  output [31:0] io_dir_req_bits_addr,
  input         io_dir_resp_bits_hit,
  input  [7:0]  io_dir_resp_bits_chosenWay,
  input         io_dir_resp_bits_isDirtyWay,
  input  [19:0] io_dir_resp_bits_tagRdVec_0,
  input  [19:0] io_dir_resp_bits_tagRdVec_1,
  input  [19:0] io_dir_resp_bits_tagRdVec_2,
  input  [19:0] io_dir_resp_bits_tagRdVec_3,
  input  [19:0] io_dir_resp_bits_tagRdVec_4,
  input  [19:0] io_dir_resp_bits_tagRdVec_5,
  input  [19:0] io_dir_resp_bits_tagRdVec_6,
  input  [19:0] io_dir_resp_bits_tagRdVec_7,
  input         io_dataBank_req_ready,
  output        io_dataBank_req_valid,
  output [7:0]  io_dataBank_req_bits_set,
  input  [31:0] io_dataBank_resp_0_0,
  input  [31:0] io_dataBank_resp_0_1,
  input  [31:0] io_dataBank_resp_0_2,
  input  [31:0] io_dataBank_resp_0_3,
  input  [31:0] io_dataBank_resp_1_0,
  input  [31:0] io_dataBank_resp_1_1,
  input  [31:0] io_dataBank_resp_1_2,
  input  [31:0] io_dataBank_resp_1_3,
  input  [31:0] io_dataBank_resp_2_0,
  input  [31:0] io_dataBank_resp_2_1,
  input  [31:0] io_dataBank_resp_2_2,
  input  [31:0] io_dataBank_resp_2_3,
  input  [31:0] io_dataBank_resp_3_0,
  input  [31:0] io_dataBank_resp_3_1,
  input  [31:0] io_dataBank_resp_3_2,
  input  [31:0] io_dataBank_resp_3_3,
  input  [31:0] io_dataBank_resp_4_0,
  input  [31:0] io_dataBank_resp_4_1,
  input  [31:0] io_dataBank_resp_4_2,
  input  [31:0] io_dataBank_resp_4_3,
  input  [31:0] io_dataBank_resp_5_0,
  input  [31:0] io_dataBank_resp_5_1,
  input  [31:0] io_dataBank_resp_5_2,
  input  [31:0] io_dataBank_resp_5_3,
  input  [31:0] io_dataBank_resp_6_0,
  input  [31:0] io_dataBank_resp_6_1,
  input  [31:0] io_dataBank_resp_6_2,
  input  [31:0] io_dataBank_resp_6_3,
  input  [31:0] io_dataBank_resp_7_0,
  input  [31:0] io_dataBank_resp_7_1,
  input  [31:0] io_dataBank_resp_7_2,
  input  [31:0] io_dataBank_resp_7_3,
  input         io_mshr_ready,
  output        io_mshr_valid,
  output [31:0] io_mshr_bits_addr,
  output        io_mshr_bits_dirInfo_hit,
  output [7:0]  io_mshr_bits_dirInfo_chosenWay,
  output        io_mshr_bits_dirInfo_isDirtyWay,
  output [19:0] io_mshr_bits_dirtyTag,
  output [31:0] io_mshr_bits_data_0,
  output [31:0] io_mshr_bits_data_1,
  output [31:0] io_mshr_bits_data_2,
  output [31:0] io_mshr_bits_data_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
`endif // RANDOMIZE_REG_INIT
  reg  s0_full; // @[LoadPipe.scala 31:26]
  wire  s0_latch = io_load_req_ready & io_load_req_valid; // @[Decoupled.scala 51:35]
  reg  s0_valid_REG; // @[LoadPipe.scala 55:25]
  reg  s0_validReg; // @[LoadPipe.scala 52:30]
  wire  _s0_valid_T_1 = io_dir_req_ready & io_dir_req_valid; // @[Decoupled.scala 51:35]
  wire  _s0_valid_T_3 = io_dataBank_req_ready & io_dataBank_req_valid; // @[Decoupled.scala 51:35]
  wire  s0_valid = (s0_valid_REG | s0_validReg) & _s0_valid_T_1 & _s0_valid_T_3; // @[LoadPipe.scala 55:71]
  reg  s1_full; // @[LoadPipe.scala 61:26]
  reg  s1_dirInfo_hit; // @[Reg.scala 19:16]
  wire  _s1_valid_T = ~s1_dirInfo_hit; // @[LoadPipe.scala 92:21]
  wire  _s1_valid_T_1 = io_mshr_ready & io_mshr_valid; // @[Decoupled.scala 51:35]
  wire  _s1_valid_T_4 = s1_dirInfo_hit & io_load_resp_valid; // @[LoadPipe.scala 93:30]
  wire  _s1_valid_T_5 = ~s1_dirInfo_hit & _s1_valid_T_1 | _s1_valid_T_4; // @[LoadPipe.scala 92:47]
  wire  s1_fire = s1_full & _s1_valid_T_5; // @[LoadPipe.scala 91:25]
  wire  s1_ready = ~s1_full | s1_fire; // @[LoadPipe.scala 75:26]
  wire  s0_fire = s0_valid & s1_ready; // @[LoadPipe.scala 33:28]
  reg [31:0] s0_reqReg_addr; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = s0_latch ? io_load_req_bits_addr : s0_reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_1 = s0_full & s0_fire ? 1'h0 : s0_full; // @[LoadPipe.scala 31:26 40:{35,45}]
  wire  _GEN_2 = s0_latch | _GEN_1; // @[LoadPipe.scala 39:{20,30}]
  wire  _GEN_3 = s0_fire ? 1'h0 : s0_validReg; // @[LoadPipe.scala 54:24 52:30 54:38]
  wire  _GEN_4 = s0_latch | _GEN_3; // @[LoadPipe.scala 53:{20,34}]
  reg [31:0] s1_rAddr; // @[Reg.scala 19:16]
  wire [3:0] s1_blockSel = 4'h1 << s1_rAddr[3:2]; // @[OneHot.scala 57:35]
  reg [31:0] s1_rdDataAll_0_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_4_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_4_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_4_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_4_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_5_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_5_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_5_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_5_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_6_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_6_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_6_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_6_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_7_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_7_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_7_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_7_3; // @[Reg.scala 19:16]
  reg [7:0] s1_dirInfo_chosenWay; // @[Reg.scala 19:16]
  reg  s1_dirInfo_isDirtyWay; // @[Reg.scala 19:16]
  wire [31:0] _s1_rdBlockData_T_8 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_9 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_10 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_11 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_12 = s1_dirInfo_chosenWay[4] ? s1_rdDataAll_4_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_13 = s1_dirInfo_chosenWay[5] ? s1_rdDataAll_5_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_14 = s1_dirInfo_chosenWay[6] ? s1_rdDataAll_6_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_15 = s1_dirInfo_chosenWay[7] ? s1_rdDataAll_7_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_16 = _s1_rdBlockData_T_8 | _s1_rdBlockData_T_9; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_17 = _s1_rdBlockData_T_16 | _s1_rdBlockData_T_10; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_18 = _s1_rdBlockData_T_17 | _s1_rdBlockData_T_11; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_19 = _s1_rdBlockData_T_18 | _s1_rdBlockData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_20 = _s1_rdBlockData_T_19 | _s1_rdBlockData_T_13; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_21 = _s1_rdBlockData_T_20 | _s1_rdBlockData_T_14; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_0 = _s1_rdBlockData_T_21 | _s1_rdBlockData_T_15; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_23 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_24 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_25 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_26 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_27 = s1_dirInfo_chosenWay[4] ? s1_rdDataAll_4_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_28 = s1_dirInfo_chosenWay[5] ? s1_rdDataAll_5_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_29 = s1_dirInfo_chosenWay[6] ? s1_rdDataAll_6_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_30 = s1_dirInfo_chosenWay[7] ? s1_rdDataAll_7_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_31 = _s1_rdBlockData_T_23 | _s1_rdBlockData_T_24; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_32 = _s1_rdBlockData_T_31 | _s1_rdBlockData_T_25; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_33 = _s1_rdBlockData_T_32 | _s1_rdBlockData_T_26; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_34 = _s1_rdBlockData_T_33 | _s1_rdBlockData_T_27; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_35 = _s1_rdBlockData_T_34 | _s1_rdBlockData_T_28; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_36 = _s1_rdBlockData_T_35 | _s1_rdBlockData_T_29; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_1 = _s1_rdBlockData_T_36 | _s1_rdBlockData_T_30; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_38 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_39 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_40 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_41 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_42 = s1_dirInfo_chosenWay[4] ? s1_rdDataAll_4_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_43 = s1_dirInfo_chosenWay[5] ? s1_rdDataAll_5_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_44 = s1_dirInfo_chosenWay[6] ? s1_rdDataAll_6_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_45 = s1_dirInfo_chosenWay[7] ? s1_rdDataAll_7_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_46 = _s1_rdBlockData_T_38 | _s1_rdBlockData_T_39; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_47 = _s1_rdBlockData_T_46 | _s1_rdBlockData_T_40; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_48 = _s1_rdBlockData_T_47 | _s1_rdBlockData_T_41; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_49 = _s1_rdBlockData_T_48 | _s1_rdBlockData_T_42; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_50 = _s1_rdBlockData_T_49 | _s1_rdBlockData_T_43; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_51 = _s1_rdBlockData_T_50 | _s1_rdBlockData_T_44; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_2 = _s1_rdBlockData_T_51 | _s1_rdBlockData_T_45; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_53 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_54 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_55 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_56 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_57 = s1_dirInfo_chosenWay[4] ? s1_rdDataAll_4_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_58 = s1_dirInfo_chosenWay[5] ? s1_rdDataAll_5_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_59 = s1_dirInfo_chosenWay[6] ? s1_rdDataAll_6_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_60 = s1_dirInfo_chosenWay[7] ? s1_rdDataAll_7_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_61 = _s1_rdBlockData_T_53 | _s1_rdBlockData_T_54; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_62 = _s1_rdBlockData_T_61 | _s1_rdBlockData_T_55; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_63 = _s1_rdBlockData_T_62 | _s1_rdBlockData_T_56; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_64 = _s1_rdBlockData_T_63 | _s1_rdBlockData_T_57; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_65 = _s1_rdBlockData_T_64 | _s1_rdBlockData_T_58; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_66 = _s1_rdBlockData_T_65 | _s1_rdBlockData_T_59; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_3 = _s1_rdBlockData_T_66 | _s1_rdBlockData_T_60; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_4 = s1_blockSel[0] ? s1_rdBlockData_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_5 = s1_blockSel[1] ? s1_rdBlockData_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_6 = s1_blockSel[2] ? s1_rdBlockData_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_7 = s1_blockSel[3] ? s1_rdBlockData_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_8 = _s1_rdData_T_4 | _s1_rdData_T_5; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_9 = _s1_rdData_T_8 | _s1_rdData_T_6; // @[Mux.scala 27:73]
  reg [19:0] s1_tagRdVec_0; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_1; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_2; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_3; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_4; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_5; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_6; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_7; // @[Reg.scala 19:16]
  wire [19:0] _s1_dirtyTag_T_8 = s1_dirInfo_chosenWay[0] ? s1_tagRdVec_0 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_9 = s1_dirInfo_chosenWay[1] ? s1_tagRdVec_1 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_10 = s1_dirInfo_chosenWay[2] ? s1_tagRdVec_2 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_11 = s1_dirInfo_chosenWay[3] ? s1_tagRdVec_3 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_12 = s1_dirInfo_chosenWay[4] ? s1_tagRdVec_4 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_13 = s1_dirInfo_chosenWay[5] ? s1_tagRdVec_5 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_14 = s1_dirInfo_chosenWay[6] ? s1_tagRdVec_6 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_15 = s1_dirInfo_chosenWay[7] ? s1_tagRdVec_7 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_16 = _s1_dirtyTag_T_8 | _s1_dirtyTag_T_9; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_17 = _s1_dirtyTag_T_16 | _s1_dirtyTag_T_10; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_18 = _s1_dirtyTag_T_17 | _s1_dirtyTag_T_11; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_19 = _s1_dirtyTag_T_18 | _s1_dirtyTag_T_12; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_20 = _s1_dirtyTag_T_19 | _s1_dirtyTag_T_13; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_21 = _s1_dirtyTag_T_20 | _s1_dirtyTag_T_14; // @[Mux.scala 27:73]
  wire  _GEN_57 = s1_full & s1_fire ? 1'h0 : s1_full; // @[LoadPipe.scala 61:26 77:{35,45}]
  wire  _GEN_58 = s0_fire | _GEN_57; // @[LoadPipe.scala 76:{20,30}]
  assign io_load_req_ready = ~s0_full; // @[LoadPipe.scala 37:26]
  assign io_load_resp_valid = s1_dirInfo_hit & s1_full; // @[LoadPipe.scala 87:36]
  assign io_load_resp_bits_data = _s1_rdData_T_9 | _s1_rdData_T_7; // @[Mux.scala 27:73]
  assign io_dir_req_valid = s0_latch | s0_full; // @[LoadPipe.scala 43:34]
  assign io_dir_req_bits_addr = s0_latch ? io_load_req_bits_addr : s0_reqReg_addr; // @[LoadPipe.scala 35:23]
  assign io_dataBank_req_valid = s0_latch | s0_full; // @[LoadPipe.scala 46:39]
  assign io_dataBank_req_bits_set = _GEN_0[11:4]; // @[Parameters.scala 50:11]
  assign io_mshr_valid = _s1_valid_T & s1_full; // @[LoadPipe.scala 79:32]
  assign io_mshr_bits_addr = s1_rAddr; // @[LoadPipe.scala 81:23]
  assign io_mshr_bits_dirInfo_hit = s1_dirInfo_hit; // @[LoadPipe.scala 84:26]
  assign io_mshr_bits_dirInfo_chosenWay = s1_dirInfo_chosenWay; // @[LoadPipe.scala 84:26]
  assign io_mshr_bits_dirInfo_isDirtyWay = s1_dirInfo_isDirtyWay; // @[LoadPipe.scala 84:26]
  assign io_mshr_bits_dirtyTag = _s1_dirtyTag_T_21 | _s1_dirtyTag_T_15; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_0 = _s1_rdBlockData_T_21 | _s1_rdBlockData_T_15; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_1 = _s1_rdBlockData_T_36 | _s1_rdBlockData_T_30; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_2 = _s1_rdBlockData_T_51 | _s1_rdBlockData_T_45; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_3 = _s1_rdBlockData_T_66 | _s1_rdBlockData_T_60; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[LoadPipe.scala 31:26]
      s0_full <= 1'h0; // @[LoadPipe.scala 31:26]
    end else begin
      s0_full <= _GEN_2;
    end
    s0_valid_REG <= io_load_req_ready & io_load_req_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[LoadPipe.scala 52:30]
      s0_validReg <= 1'h0; // @[LoadPipe.scala 52:30]
    end else begin
      s0_validReg <= _GEN_4;
    end
    if (reset) begin // @[LoadPipe.scala 61:26]
      s1_full <= 1'h0; // @[LoadPipe.scala 61:26]
    end else begin
      s1_full <= _GEN_58;
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_hit <= io_dir_resp_bits_hit; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_addr <= io_load_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      if (s0_latch) begin // @[Reg.scala 20:18]
        s1_rAddr <= io_load_req_bits_addr; // @[Reg.scala 20:22]
      end else begin
        s1_rAddr <= s0_reqReg_addr; // @[Reg.scala 19:16]
      end
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_0 <= io_dataBank_resp_0_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_1 <= io_dataBank_resp_0_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_2 <= io_dataBank_resp_0_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_3 <= io_dataBank_resp_0_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_0 <= io_dataBank_resp_1_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_1 <= io_dataBank_resp_1_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_2 <= io_dataBank_resp_1_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_3 <= io_dataBank_resp_1_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_0 <= io_dataBank_resp_2_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_1 <= io_dataBank_resp_2_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_2 <= io_dataBank_resp_2_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_3 <= io_dataBank_resp_2_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_0 <= io_dataBank_resp_3_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_1 <= io_dataBank_resp_3_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_2 <= io_dataBank_resp_3_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_3 <= io_dataBank_resp_3_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_4_0 <= io_dataBank_resp_4_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_4_1 <= io_dataBank_resp_4_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_4_2 <= io_dataBank_resp_4_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_4_3 <= io_dataBank_resp_4_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_5_0 <= io_dataBank_resp_5_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_5_1 <= io_dataBank_resp_5_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_5_2 <= io_dataBank_resp_5_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_5_3 <= io_dataBank_resp_5_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_6_0 <= io_dataBank_resp_6_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_6_1 <= io_dataBank_resp_6_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_6_2 <= io_dataBank_resp_6_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_6_3 <= io_dataBank_resp_6_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_7_0 <= io_dataBank_resp_7_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_7_1 <= io_dataBank_resp_7_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_7_2 <= io_dataBank_resp_7_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_7_3 <= io_dataBank_resp_7_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_chosenWay <= io_dir_resp_bits_chosenWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_isDirtyWay <= io_dir_resp_bits_isDirtyWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_0 <= io_dir_resp_bits_tagRdVec_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_1 <= io_dir_resp_bits_tagRdVec_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_2 <= io_dir_resp_bits_tagRdVec_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_3 <= io_dir_resp_bits_tagRdVec_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_4 <= io_dir_resp_bits_tagRdVec_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_5 <= io_dir_resp_bits_tagRdVec_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_6 <= io_dir_resp_bits_tagRdVec_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_7 <= io_dir_resp_bits_tagRdVec_7; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s0_valid_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s0_validReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s1_full = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s1_dirInfo_hit = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s0_reqReg_addr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  s1_rAddr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  s1_rdDataAll_0_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  s1_rdDataAll_0_1 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  s1_rdDataAll_0_2 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  s1_rdDataAll_0_3 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  s1_rdDataAll_1_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  s1_rdDataAll_1_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  s1_rdDataAll_1_2 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  s1_rdDataAll_1_3 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  s1_rdDataAll_2_0 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  s1_rdDataAll_2_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  s1_rdDataAll_2_2 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  s1_rdDataAll_2_3 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  s1_rdDataAll_3_0 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  s1_rdDataAll_3_1 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  s1_rdDataAll_3_2 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  s1_rdDataAll_3_3 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  s1_rdDataAll_4_0 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  s1_rdDataAll_4_1 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  s1_rdDataAll_4_2 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  s1_rdDataAll_4_3 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  s1_rdDataAll_5_0 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  s1_rdDataAll_5_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  s1_rdDataAll_5_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  s1_rdDataAll_5_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  s1_rdDataAll_6_0 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  s1_rdDataAll_6_1 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  s1_rdDataAll_6_2 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  s1_rdDataAll_6_3 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  s1_rdDataAll_7_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  s1_rdDataAll_7_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  s1_rdDataAll_7_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  s1_rdDataAll_7_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  s1_dirInfo_chosenWay = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  s1_dirInfo_isDirtyWay = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  s1_tagRdVec_0 = _RAND_41[19:0];
  _RAND_42 = {1{`RANDOM}};
  s1_tagRdVec_1 = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  s1_tagRdVec_2 = _RAND_43[19:0];
  _RAND_44 = {1{`RANDOM}};
  s1_tagRdVec_3 = _RAND_44[19:0];
  _RAND_45 = {1{`RANDOM}};
  s1_tagRdVec_4 = _RAND_45[19:0];
  _RAND_46 = {1{`RANDOM}};
  s1_tagRdVec_5 = _RAND_46[19:0];
  _RAND_47 = {1{`RANDOM}};
  s1_tagRdVec_6 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  s1_tagRdVec_7 = _RAND_48[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StorePipe(
  input         clock,
  input         reset,
  output        io_store_req_ready,
  input         io_store_req_valid,
  input  [31:0] io_store_req_bits_addr,
  input  [31:0] io_store_req_bits_data,
  input  [3:0]  io_store_req_bits_mask,
  output        io_store_resp_valid,
  output        io_dir_read_req_valid,
  output [31:0] io_dir_read_req_bits_addr,
  input         io_dir_read_resp_bits_hit,
  input  [7:0]  io_dir_read_resp_bits_chosenWay,
  input         io_dir_read_resp_bits_isDirtyWay,
  input  [19:0] io_dir_read_resp_bits_tagRdVec_0,
  input  [19:0] io_dir_read_resp_bits_tagRdVec_1,
  input  [19:0] io_dir_read_resp_bits_tagRdVec_2,
  input  [19:0] io_dir_read_resp_bits_tagRdVec_3,
  input  [19:0] io_dir_read_resp_bits_tagRdVec_4,
  input  [19:0] io_dir_read_resp_bits_tagRdVec_5,
  input  [19:0] io_dir_read_resp_bits_tagRdVec_6,
  input  [19:0] io_dir_read_resp_bits_tagRdVec_7,
  output        io_dir_write_req_valid,
  output [31:0] io_dir_write_req_bits_addr,
  output [7:0]  io_dir_write_req_bits_way,
  output        io_dataBank_read_req_valid,
  output [7:0]  io_dataBank_read_req_bits_set,
  input  [31:0] io_dataBank_read_resp_0_0,
  input  [31:0] io_dataBank_read_resp_0_1,
  input  [31:0] io_dataBank_read_resp_0_2,
  input  [31:0] io_dataBank_read_resp_0_3,
  input  [31:0] io_dataBank_read_resp_1_0,
  input  [31:0] io_dataBank_read_resp_1_1,
  input  [31:0] io_dataBank_read_resp_1_2,
  input  [31:0] io_dataBank_read_resp_1_3,
  input  [31:0] io_dataBank_read_resp_2_0,
  input  [31:0] io_dataBank_read_resp_2_1,
  input  [31:0] io_dataBank_read_resp_2_2,
  input  [31:0] io_dataBank_read_resp_2_3,
  input  [31:0] io_dataBank_read_resp_3_0,
  input  [31:0] io_dataBank_read_resp_3_1,
  input  [31:0] io_dataBank_read_resp_3_2,
  input  [31:0] io_dataBank_read_resp_3_3,
  input  [31:0] io_dataBank_read_resp_4_0,
  input  [31:0] io_dataBank_read_resp_4_1,
  input  [31:0] io_dataBank_read_resp_4_2,
  input  [31:0] io_dataBank_read_resp_4_3,
  input  [31:0] io_dataBank_read_resp_5_0,
  input  [31:0] io_dataBank_read_resp_5_1,
  input  [31:0] io_dataBank_read_resp_5_2,
  input  [31:0] io_dataBank_read_resp_5_3,
  input  [31:0] io_dataBank_read_resp_6_0,
  input  [31:0] io_dataBank_read_resp_6_1,
  input  [31:0] io_dataBank_read_resp_6_2,
  input  [31:0] io_dataBank_read_resp_6_3,
  input  [31:0] io_dataBank_read_resp_7_0,
  input  [31:0] io_dataBank_read_resp_7_1,
  input  [31:0] io_dataBank_read_resp_7_2,
  input  [31:0] io_dataBank_read_resp_7_3,
  output        io_dataBank_write_req_valid,
  output [7:0]  io_dataBank_write_req_bits_set,
  output [31:0] io_dataBank_write_req_bits_data_0,
  output [31:0] io_dataBank_write_req_bits_data_1,
  output [31:0] io_dataBank_write_req_bits_data_2,
  output [31:0] io_dataBank_write_req_bits_data_3,
  output [3:0]  io_dataBank_write_req_bits_blockMask,
  output [7:0]  io_dataBank_write_req_bits_way,
  input         io_mshr_ready,
  output        io_mshr_valid,
  output [31:0] io_mshr_bits_addr,
  output        io_mshr_bits_dirInfo_hit,
  output [7:0]  io_mshr_bits_dirInfo_chosenWay,
  output        io_mshr_bits_dirInfo_isDirtyWay,
  output [19:0] io_mshr_bits_dirtyTag,
  output [31:0] io_mshr_bits_data_0,
  output [31:0] io_mshr_bits_data_1,
  output [31:0] io_mshr_bits_data_2,
  output [31:0] io_mshr_bits_data_3,
  output [31:0] io_mshr_bits_storeData,
  output [3:0]  io_mshr_bits_storeMask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
`endif // RANDOMIZE_REG_INIT
  reg  s0_full; // @[StorePipe.scala 30:26]
  wire  s0_latch = io_store_req_ready & io_store_req_valid; // @[Decoupled.scala 51:35]
  reg  s0_valid_REG; // @[StorePipe.scala 56:25]
  reg  s0_validReg; // @[StorePipe.scala 53:30]
  wire  s0_valid = (s0_valid_REG | s0_validReg) & io_dir_read_req_valid & io_dataBank_read_req_valid; // @[StorePipe.scala 56:77]
  reg  s1_full; // @[StorePipe.scala 63:26]
  reg  s1_dirInfo_hit; // @[Reg.scala 19:16]
  wire  _s1_valid_T = ~s1_dirInfo_hit; // @[StorePipe.scala 114:21]
  wire  _s1_valid_T_1 = io_mshr_ready & io_mshr_valid; // @[Decoupled.scala 51:35]
  wire  _s1_valid_T_6 = s1_dirInfo_hit & io_dataBank_write_req_valid & io_dir_write_req_valid; // @[StorePipe.scala 115:60]
  wire  _s1_valid_T_7 = ~s1_dirInfo_hit & _s1_valid_T_1 | _s1_valid_T_6; // @[StorePipe.scala 114:47]
  wire  s1_valid = s1_full & _s1_valid_T_7; // @[StorePipe.scala 113:25]
  reg  s2_full; // @[StorePipe.scala 121:26]
  reg  s2_isHit; // @[Reg.scala 19:16]
  wire  s2_fire = io_store_resp_valid & s2_full & s2_isHit | ~s2_isHit; // @[StorePipe.scala 133:59]
  wire  s2_ready = ~s2_full | s2_fire; // @[StorePipe.scala 126:26]
  wire  s1_fire = s1_valid & s2_ready; // @[StorePipe.scala 65:28]
  wire  s1_ready = ~s1_full | s1_fire; // @[StorePipe.scala 80:26]
  wire  s0_fire = s0_valid & s1_ready; // @[StorePipe.scala 32:28]
  reg [31:0] s0_reqReg_addr; // @[Reg.scala 19:16]
  reg [31:0] s0_reqReg_data; // @[Reg.scala 19:16]
  reg [3:0] s0_reqReg_mask; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = s0_latch ? io_store_req_bits_addr : s0_reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_3 = s0_full & s0_fire ? 1'h0 : s0_full; // @[StorePipe.scala 30:26 40:{35,45}]
  wire  _GEN_4 = s0_latch | _GEN_3; // @[StorePipe.scala 39:{20,30}]
  wire  _GEN_5 = s0_fire ? 1'h0 : s0_validReg; // @[StorePipe.scala 55:24 53:30 55:38]
  wire  _GEN_6 = s0_latch | _GEN_5; // @[StorePipe.scala 54:{20,34}]
  reg [31:0] s1_reqReg_addr; // @[Reg.scala 19:16]
  reg [31:0] s1_reqReg_data; // @[Reg.scala 19:16]
  reg [3:0] s1_reqReg_mask; // @[Reg.scala 19:16]
  wire [3:0] s1_dataBlockSelOH = 4'h1 << s1_reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  reg [31:0] s1_rdDataAll_0_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_0_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_1_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_2_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_3_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_4_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_4_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_4_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_4_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_5_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_5_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_5_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_5_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_6_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_6_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_6_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_6_3; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_7_0; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_7_1; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_7_2; // @[Reg.scala 19:16]
  reg [31:0] s1_rdDataAll_7_3; // @[Reg.scala 19:16]
  reg [7:0] s1_dirInfo_chosenWay; // @[Reg.scala 19:16]
  reg  s1_dirInfo_isDirtyWay; // @[Reg.scala 19:16]
  wire [31:0] _s1_rdBlockData_T_8 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_9 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_10 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_11 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_12 = s1_dirInfo_chosenWay[4] ? s1_rdDataAll_4_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_13 = s1_dirInfo_chosenWay[5] ? s1_rdDataAll_5_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_14 = s1_dirInfo_chosenWay[6] ? s1_rdDataAll_6_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_15 = s1_dirInfo_chosenWay[7] ? s1_rdDataAll_7_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_16 = _s1_rdBlockData_T_8 | _s1_rdBlockData_T_9; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_17 = _s1_rdBlockData_T_16 | _s1_rdBlockData_T_10; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_18 = _s1_rdBlockData_T_17 | _s1_rdBlockData_T_11; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_19 = _s1_rdBlockData_T_18 | _s1_rdBlockData_T_12; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_20 = _s1_rdBlockData_T_19 | _s1_rdBlockData_T_13; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_21 = _s1_rdBlockData_T_20 | _s1_rdBlockData_T_14; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_0 = _s1_rdBlockData_T_21 | _s1_rdBlockData_T_15; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_23 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_24 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_25 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_26 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_27 = s1_dirInfo_chosenWay[4] ? s1_rdDataAll_4_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_28 = s1_dirInfo_chosenWay[5] ? s1_rdDataAll_5_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_29 = s1_dirInfo_chosenWay[6] ? s1_rdDataAll_6_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_30 = s1_dirInfo_chosenWay[7] ? s1_rdDataAll_7_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_31 = _s1_rdBlockData_T_23 | _s1_rdBlockData_T_24; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_32 = _s1_rdBlockData_T_31 | _s1_rdBlockData_T_25; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_33 = _s1_rdBlockData_T_32 | _s1_rdBlockData_T_26; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_34 = _s1_rdBlockData_T_33 | _s1_rdBlockData_T_27; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_35 = _s1_rdBlockData_T_34 | _s1_rdBlockData_T_28; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_36 = _s1_rdBlockData_T_35 | _s1_rdBlockData_T_29; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_1 = _s1_rdBlockData_T_36 | _s1_rdBlockData_T_30; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_38 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_39 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_40 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_41 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_42 = s1_dirInfo_chosenWay[4] ? s1_rdDataAll_4_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_43 = s1_dirInfo_chosenWay[5] ? s1_rdDataAll_5_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_44 = s1_dirInfo_chosenWay[6] ? s1_rdDataAll_6_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_45 = s1_dirInfo_chosenWay[7] ? s1_rdDataAll_7_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_46 = _s1_rdBlockData_T_38 | _s1_rdBlockData_T_39; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_47 = _s1_rdBlockData_T_46 | _s1_rdBlockData_T_40; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_48 = _s1_rdBlockData_T_47 | _s1_rdBlockData_T_41; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_49 = _s1_rdBlockData_T_48 | _s1_rdBlockData_T_42; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_50 = _s1_rdBlockData_T_49 | _s1_rdBlockData_T_43; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_51 = _s1_rdBlockData_T_50 | _s1_rdBlockData_T_44; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_2 = _s1_rdBlockData_T_51 | _s1_rdBlockData_T_45; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_53 = s1_dirInfo_chosenWay[0] ? s1_rdDataAll_0_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_54 = s1_dirInfo_chosenWay[1] ? s1_rdDataAll_1_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_55 = s1_dirInfo_chosenWay[2] ? s1_rdDataAll_2_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_56 = s1_dirInfo_chosenWay[3] ? s1_rdDataAll_3_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_57 = s1_dirInfo_chosenWay[4] ? s1_rdDataAll_4_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_58 = s1_dirInfo_chosenWay[5] ? s1_rdDataAll_5_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_59 = s1_dirInfo_chosenWay[6] ? s1_rdDataAll_6_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_60 = s1_dirInfo_chosenWay[7] ? s1_rdDataAll_7_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_61 = _s1_rdBlockData_T_53 | _s1_rdBlockData_T_54; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_62 = _s1_rdBlockData_T_61 | _s1_rdBlockData_T_55; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_63 = _s1_rdBlockData_T_62 | _s1_rdBlockData_T_56; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_64 = _s1_rdBlockData_T_63 | _s1_rdBlockData_T_57; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_65 = _s1_rdBlockData_T_64 | _s1_rdBlockData_T_58; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdBlockData_T_66 = _s1_rdBlockData_T_65 | _s1_rdBlockData_T_59; // @[Mux.scala 27:73]
  wire [31:0] s1_rdBlockData_3 = _s1_rdBlockData_T_66 | _s1_rdBlockData_T_60; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_4 = s1_dataBlockSelOH[0] ? s1_rdBlockData_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_5 = s1_dataBlockSelOH[1] ? s1_rdBlockData_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_6 = s1_dataBlockSelOH[2] ? s1_rdBlockData_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_7 = s1_dataBlockSelOH[3] ? s1_rdBlockData_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_8 = _s1_rdData_T_4 | _s1_rdData_T_5; // @[Mux.scala 27:73]
  wire [31:0] _s1_rdData_T_9 = _s1_rdData_T_8 | _s1_rdData_T_6; // @[Mux.scala 27:73]
  wire [31:0] s1_rdData = _s1_rdData_T_9 | _s1_rdData_T_7; // @[Mux.scala 27:73]
  reg [19:0] s1_tagRdVec_0; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_1; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_2; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_3; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_4; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_5; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_6; // @[Reg.scala 19:16]
  reg [19:0] s1_tagRdVec_7; // @[Reg.scala 19:16]
  wire [19:0] _s1_dirtyTag_T_8 = s1_dirInfo_chosenWay[0] ? s1_tagRdVec_0 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_9 = s1_dirInfo_chosenWay[1] ? s1_tagRdVec_1 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_10 = s1_dirInfo_chosenWay[2] ? s1_tagRdVec_2 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_11 = s1_dirInfo_chosenWay[3] ? s1_tagRdVec_3 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_12 = s1_dirInfo_chosenWay[4] ? s1_tagRdVec_4 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_13 = s1_dirInfo_chosenWay[5] ? s1_tagRdVec_5 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_14 = s1_dirInfo_chosenWay[6] ? s1_tagRdVec_6 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_15 = s1_dirInfo_chosenWay[7] ? s1_tagRdVec_7 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_16 = _s1_dirtyTag_T_8 | _s1_dirtyTag_T_9; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_17 = _s1_dirtyTag_T_16 | _s1_dirtyTag_T_10; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_18 = _s1_dirtyTag_T_17 | _s1_dirtyTag_T_11; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_19 = _s1_dirtyTag_T_18 | _s1_dirtyTag_T_12; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_20 = _s1_dirtyTag_T_19 | _s1_dirtyTag_T_13; // @[Mux.scala 27:73]
  wire [19:0] _s1_dirtyTag_T_21 = _s1_dirtyTag_T_20 | _s1_dirtyTag_T_14; // @[Mux.scala 27:73]
  wire  _GEN_61 = s1_full & s1_fire ? 1'h0 : s1_full; // @[StorePipe.scala 63:26 82:{35,45}]
  wire  _GEN_62 = s0_fire | _GEN_61; // @[StorePipe.scala 81:{20,30}]
  wire [1:0] hi = s1_dataBlockSelOH[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo = s1_dataBlockSelOH[1:0]; // @[OneHot.scala 31:18]
  wire  _T_2 = |hi; // @[OneHot.scala 32:14]
  wire [1:0] _T_3 = hi | lo; // @[OneHot.scala 32:28]
  wire [1:0] _T_5 = {_T_2,_T_3[1]}; // @[Cat.scala 33:92]
  wire [7:0] _tempWrData_tempMask_T_5 = s1_reqReg_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_7 = s1_reqReg_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_9 = s1_reqReg_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_11 = s1_reqReg_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [31:0] tempWrData_tempMask = {_tempWrData_tempMask_T_11,_tempWrData_tempMask_T_9,_tempWrData_tempMask_T_7,
    _tempWrData_tempMask_T_5}; // @[Cat.scala 33:92]
  wire [31:0] _tempWrData_T = ~tempWrData_tempMask; // @[Parameters.scala 67:8]
  wire [31:0] _tempWrData_T_1 = _tempWrData_T & s1_rdData; // @[Parameters.scala 67:18]
  wire [31:0] _tempWrData_T_2 = tempWrData_tempMask & s1_reqReg_data; // @[Parameters.scala 67:41]
  wire [31:0] _tempWrData_T_3 = _tempWrData_T_1 | _tempWrData_T_2; // @[Parameters.scala 67:29]
  wire  _GEN_68 = s2_full & s2_fire ? 1'h0 : s2_full; // @[StorePipe.scala 121:26 128:{35,45}]
  wire  _GEN_69 = s1_fire | _GEN_68; // @[StorePipe.scala 127:{20,30}]
  assign io_store_req_ready = ~s0_full; // @[StorePipe.scala 38:27]
  assign io_store_resp_valid = s2_isHit & s2_full; // @[StorePipe.scala 130:37]
  assign io_dir_read_req_valid = s0_latch | s0_full; // @[StorePipe.scala 43:39]
  assign io_dir_read_req_bits_addr = s0_latch ? io_store_req_bits_addr : s0_reqReg_addr; // @[StorePipe.scala 34:23]
  assign io_dir_write_req_valid = s1_dirInfo_hit & s1_full; // @[StorePipe.scala 94:40]
  assign io_dir_write_req_bits_addr = s1_reqReg_addr; // @[StorePipe.scala 96:32]
  assign io_dir_write_req_bits_way = s1_dirInfo_chosenWay; // @[StorePipe.scala 101:31]
  assign io_dataBank_read_req_valid = s0_latch | s0_full; // @[StorePipe.scala 46:44]
  assign io_dataBank_read_req_bits_set = _GEN_0[11:4]; // @[Parameters.scala 50:11]
  assign io_dataBank_write_req_valid = s1_dirInfo_hit & s1_full; // @[StorePipe.scala 103:45]
  assign io_dataBank_write_req_bits_set = s1_reqReg_addr[11:4]; // @[Parameters.scala 50:11]
  assign io_dataBank_write_req_bits_data_0 = 2'h0 == _T_5 ? _tempWrData_T_3 : 32'h0; // @[StorePipe.scala 108:30 109:{45,45}]
  assign io_dataBank_write_req_bits_data_1 = 2'h1 == _T_5 ? _tempWrData_T_3 : 32'h0; // @[StorePipe.scala 108:30 109:{45,45}]
  assign io_dataBank_write_req_bits_data_2 = 2'h2 == _T_5 ? _tempWrData_T_3 : 32'h0; // @[StorePipe.scala 108:30 109:{45,45}]
  assign io_dataBank_write_req_bits_data_3 = 2'h3 == _T_5 ? _tempWrData_T_3 : 32'h0; // @[StorePipe.scala 108:30 109:{45,45}]
  assign io_dataBank_write_req_bits_blockMask = 4'h1 << s1_reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  assign io_dataBank_write_req_bits_way = s1_dirInfo_chosenWay; // @[StorePipe.scala 107:36]
  assign io_mshr_valid = _s1_valid_T & s1_full; // @[StorePipe.scala 84:32]
  assign io_mshr_bits_addr = s1_reqReg_addr; // @[StorePipe.scala 86:23]
  assign io_mshr_bits_dirInfo_hit = s1_dirInfo_hit; // @[StorePipe.scala 87:26]
  assign io_mshr_bits_dirInfo_chosenWay = s1_dirInfo_chosenWay; // @[StorePipe.scala 87:26]
  assign io_mshr_bits_dirInfo_isDirtyWay = s1_dirInfo_isDirtyWay; // @[StorePipe.scala 87:26]
  assign io_mshr_bits_dirtyTag = _s1_dirtyTag_T_21 | _s1_dirtyTag_T_15; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_0 = _s1_rdBlockData_T_21 | _s1_rdBlockData_T_15; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_1 = _s1_rdBlockData_T_36 | _s1_rdBlockData_T_30; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_2 = _s1_rdBlockData_T_51 | _s1_rdBlockData_T_45; // @[Mux.scala 27:73]
  assign io_mshr_bits_data_3 = _s1_rdBlockData_T_66 | _s1_rdBlockData_T_60; // @[Mux.scala 27:73]
  assign io_mshr_bits_storeData = s1_reqReg_data; // @[StorePipe.scala 91:28]
  assign io_mshr_bits_storeMask = s1_reqReg_mask; // @[StorePipe.scala 92:28]
  always @(posedge clock) begin
    if (reset) begin // @[StorePipe.scala 30:26]
      s0_full <= 1'h0; // @[StorePipe.scala 30:26]
    end else begin
      s0_full <= _GEN_4;
    end
    s0_valid_REG <= io_store_req_ready & io_store_req_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[StorePipe.scala 53:30]
      s0_validReg <= 1'h0; // @[StorePipe.scala 53:30]
    end else begin
      s0_validReg <= _GEN_6;
    end
    if (reset) begin // @[StorePipe.scala 63:26]
      s1_full <= 1'h0; // @[StorePipe.scala 63:26]
    end else begin
      s1_full <= _GEN_62;
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_hit <= io_dir_read_resp_bits_hit; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[StorePipe.scala 121:26]
      s2_full <= 1'h0; // @[StorePipe.scala 121:26]
    end else begin
      s2_full <= _GEN_69;
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_isHit <= s1_dirInfo_hit; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_addr <= io_store_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_data <= io_store_req_bits_data; // @[Reg.scala 20:22]
    end
    if (s0_latch) begin // @[Reg.scala 20:18]
      s0_reqReg_mask <= io_store_req_bits_mask; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_reqReg_addr <= s0_reqReg_addr; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_reqReg_data <= s0_reqReg_data; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_reqReg_mask <= s0_reqReg_mask; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_0 <= io_dataBank_read_resp_0_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_1 <= io_dataBank_read_resp_0_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_2 <= io_dataBank_read_resp_0_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_0_3 <= io_dataBank_read_resp_0_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_0 <= io_dataBank_read_resp_1_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_1 <= io_dataBank_read_resp_1_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_2 <= io_dataBank_read_resp_1_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_1_3 <= io_dataBank_read_resp_1_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_0 <= io_dataBank_read_resp_2_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_1 <= io_dataBank_read_resp_2_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_2 <= io_dataBank_read_resp_2_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_2_3 <= io_dataBank_read_resp_2_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_0 <= io_dataBank_read_resp_3_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_1 <= io_dataBank_read_resp_3_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_2 <= io_dataBank_read_resp_3_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_3_3 <= io_dataBank_read_resp_3_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_4_0 <= io_dataBank_read_resp_4_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_4_1 <= io_dataBank_read_resp_4_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_4_2 <= io_dataBank_read_resp_4_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_4_3 <= io_dataBank_read_resp_4_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_5_0 <= io_dataBank_read_resp_5_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_5_1 <= io_dataBank_read_resp_5_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_5_2 <= io_dataBank_read_resp_5_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_5_3 <= io_dataBank_read_resp_5_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_6_0 <= io_dataBank_read_resp_6_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_6_1 <= io_dataBank_read_resp_6_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_6_2 <= io_dataBank_read_resp_6_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_6_3 <= io_dataBank_read_resp_6_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_7_0 <= io_dataBank_read_resp_7_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_7_1 <= io_dataBank_read_resp_7_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_7_2 <= io_dataBank_read_resp_7_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_rdDataAll_7_3 <= io_dataBank_read_resp_7_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_chosenWay <= io_dir_read_resp_bits_chosenWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_dirInfo_isDirtyWay <= io_dir_read_resp_bits_isDirtyWay; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_0 <= io_dir_read_resp_bits_tagRdVec_0; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_1 <= io_dir_read_resp_bits_tagRdVec_1; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_2 <= io_dir_read_resp_bits_tagRdVec_2; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_3 <= io_dir_read_resp_bits_tagRdVec_3; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_4 <= io_dir_read_resp_bits_tagRdVec_4; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_5 <= io_dir_read_resp_bits_tagRdVec_5; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_6 <= io_dir_read_resp_bits_tagRdVec_6; // @[Reg.scala 20:22]
    end
    if (s0_fire) begin // @[Reg.scala 20:18]
      s1_tagRdVec_7 <= io_dir_read_resp_bits_tagRdVec_7; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s0_valid_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s0_validReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s1_full = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s1_dirInfo_hit = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s2_full = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s2_isHit = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s0_reqReg_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  s0_reqReg_data = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  s0_reqReg_mask = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  s1_reqReg_addr = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  s1_reqReg_data = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  s1_reqReg_mask = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  s1_rdDataAll_0_0 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  s1_rdDataAll_0_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  s1_rdDataAll_0_2 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  s1_rdDataAll_0_3 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  s1_rdDataAll_1_0 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  s1_rdDataAll_1_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  s1_rdDataAll_1_2 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  s1_rdDataAll_1_3 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  s1_rdDataAll_2_0 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  s1_rdDataAll_2_1 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  s1_rdDataAll_2_2 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  s1_rdDataAll_2_3 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  s1_rdDataAll_3_0 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  s1_rdDataAll_3_1 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  s1_rdDataAll_3_2 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  s1_rdDataAll_3_3 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  s1_rdDataAll_4_0 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  s1_rdDataAll_4_1 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  s1_rdDataAll_4_2 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  s1_rdDataAll_4_3 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  s1_rdDataAll_5_0 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  s1_rdDataAll_5_1 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  s1_rdDataAll_5_2 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  s1_rdDataAll_5_3 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  s1_rdDataAll_6_0 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  s1_rdDataAll_6_1 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  s1_rdDataAll_6_2 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  s1_rdDataAll_6_3 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  s1_rdDataAll_7_0 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  s1_rdDataAll_7_1 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  s1_rdDataAll_7_2 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  s1_rdDataAll_7_3 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  s1_dirInfo_chosenWay = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  s1_dirInfo_isDirtyWay = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  s1_tagRdVec_0 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  s1_tagRdVec_1 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  s1_tagRdVec_2 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  s1_tagRdVec_3 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  s1_tagRdVec_4 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  s1_tagRdVec_5 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  s1_tagRdVec_6 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  s1_tagRdVec_7 = _RAND_54[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MSHR(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [31:0] io_req_bits_addr,
  input         io_req_bits_dirInfo_hit,
  input  [7:0]  io_req_bits_dirInfo_chosenWay,
  input         io_req_bits_dirInfo_isDirtyWay,
  input  [19:0] io_req_bits_dirtyTag,
  input  [31:0] io_req_bits_data_0,
  input  [31:0] io_req_bits_data_1,
  input  [31:0] io_req_bits_data_2,
  input  [31:0] io_req_bits_data_3,
  input         io_req_bits_isStore,
  input  [31:0] io_req_bits_storeData,
  input  [3:0]  io_req_bits_storeMask,
  input         io_resp_load_ready,
  output        io_resp_load_valid,
  output [31:0] io_resp_load_bits_data,
  input         io_resp_store_ready,
  output        io_resp_store_valid,
  output        io_tasks_refill_req_valid,
  output [31:0] io_tasks_refill_req_bits_addr,
  output [7:0]  io_tasks_refill_req_bits_chosenWay,
  output        io_tasks_refill_resp_ready,
  input         io_tasks_refill_resp_valid,
  input  [31:0] io_tasks_refill_resp_bits_data,
  output        io_tasks_writeback_req_valid,
  output [31:0] io_tasks_writeback_req_bits_addr,
  output [19:0] io_tasks_writeback_req_bits_dirtyTag,
  output [31:0] io_tasks_writeback_req_bits_data_0,
  output [31:0] io_tasks_writeback_req_bits_data_1,
  output [31:0] io_tasks_writeback_req_bits_data_2,
  output [31:0] io_tasks_writeback_req_bits_data_3,
  output        io_tasks_writeback_resp_ready,
  input         io_tasks_writeback_resp_valid,
  input         io_dirWrite_req_ready,
  output        io_dirWrite_req_valid,
  output [31:0] io_dirWrite_req_bits_addr,
  output [7:0]  io_dirWrite_req_bits_way,
  input         io_dataWrite_req_ready,
  output        io_dataWrite_req_valid,
  output [7:0]  io_dataWrite_req_bits_set,
  output [31:0] io_dataWrite_req_bits_data_0,
  output [31:0] io_dataWrite_req_bits_data_1,
  output [31:0] io_dataWrite_req_bits_data_2,
  output [31:0] io_dataWrite_req_bits_data_3,
  output [3:0]  io_dataWrite_req_bits_blockMask,
  output [7:0]  io_dataWrite_req_bits_way
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] reqReg_addr; // @[Reg.scala 19:16]
  reg [7:0] reqReg_dirInfo_chosenWay; // @[Reg.scala 19:16]
  reg [19:0] reqReg_dirtyTag; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_0; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_1; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_2; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_3; // @[Reg.scala 19:16]
  reg  reqReg_isStore; // @[Reg.scala 19:16]
  reg [31:0] reqReg_storeData; // @[Reg.scala 19:16]
  reg [3:0] reqReg_storeMask; // @[Reg.scala 19:16]
  wire  _GEN_17 = _reqReg_T ? io_req_bits_isStore : reqReg_isStore; // @[Reg.scala 19:16 20:{18,22}]
  reg [2:0] state; // @[MSHR.scala 64:24]
  wire  _io_busy_T = state == 3'h0; // @[MSHR.scala 67:22]
  wire [1:0] _GEN_21 = io_req_bits_dirInfo_isDirtyWay ? 2'h1 : 2'h2; // @[MSHR.scala 74:50 75:27 77:27]
  wire [1:0] _GEN_22 = _reqReg_T ? _GEN_21 : 2'h0; // @[MSHR.scala 72:19 73:27]
  wire [1:0] _GEN_23 = _io_busy_T ? _GEN_22 : 2'h0; // @[MSHR.scala 71:27 65:29]
  wire  _T_2 = state == 3'h1; // @[MSHR.scala 83:16]
  wire  _T_3 = io_tasks_writeback_resp_ready & io_tasks_writeback_resp_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_24 = _T_3 ? 2'h2 : 2'h1; // @[MSHR.scala 84:19 85:44 86:23]
  wire [1:0] _GEN_25 = state == 3'h1 ? _GEN_24 : _GEN_23; // @[MSHR.scala 83:32]
  wire  _T_4 = state == 3'h2; // @[MSHR.scala 91:16]
  wire  _T_5 = io_tasks_refill_resp_ready & io_tasks_refill_resp_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_26 = _T_5 ? 3'h4 : 3'h2; // @[MSHR.scala 92:19 95:47 96:23]
  wire [2:0] _GEN_27 = _T_5 & _GEN_17 ? 3'h3 : _GEN_26; // @[MSHR.scala 93:56 94:23]
  wire  _T_8 = io_resp_load_ready & io_resp_load_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_28 = _T_8 ? 3'h0 : _GEN_27; // @[MSHR.scala 100:23 99:33]
  wire  _T_9 = state == 3'h3; // @[MSHR.scala 105:16]
  wire  _T_10 = io_dirWrite_req_ready & io_dirWrite_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_11 = io_dataWrite_req_ready & io_dataWrite_req_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_30 = _T_10 & _T_11 ? 3'h4 : 3'h3; // @[MSHR.scala 106:19 107:61 108:23]
  wire  _T_13 = io_resp_store_ready & io_resp_store_valid; // @[Decoupled.scala 51:35]
  wire  _T_14 = state == 3'h4; // @[MSHR.scala 117:16]
  wire  _willRefill_T_1 = ~io_req_bits_dirInfo_hit; // @[MSHR.scala 126:63]
  wire  willRefill = ~io_req_bits_dirInfo_isDirtyWay & ~io_req_bits_dirInfo_hit & _reqReg_T; // @[MSHR.scala 126:88]
  wire  willWriteback = io_req_bits_dirInfo_isDirtyWay & _willRefill_T_1 & _reqReg_T; // @[MSHR.scala 127:87]
  wire  willWriteStore = _T_4 & _GEN_17 & _T_5; // @[MSHR.scala 128:61]
  wire  _willRespLoad_T_1 = ~_GEN_17; // @[MSHR.scala 129:49]
  wire  willRespLoad = _T_4 & ~_GEN_17 & _T_5; // @[MSHR.scala 129:62]
  wire  willRespStore = _T_9 & _T_10 & _T_11; // @[MSHR.scala 130:73]
  wire [3:0] _io_dataWrite_req_bits_blockMask_T_1 = 4'h1 << reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  reg [31:0] oldData_r; // @[Reg.scala 19:16]
  wire [31:0] _GEN_35 = _T_5 ? io_tasks_refill_resp_bits_data : oldData_r; // @[Reg.scala 19:16 20:{18,22}]
  wire [1:0] hi = _io_dataWrite_req_bits_blockMask_T_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo = _io_dataWrite_req_bits_blockMask_T_1[1:0]; // @[OneHot.scala 31:18]
  wire  _T_20 = |hi; // @[OneHot.scala 32:14]
  wire [1:0] _T_21 = hi | lo; // @[OneHot.scala 32:28]
  wire [1:0] _T_23 = {_T_20,_T_21[1]}; // @[Cat.scala 33:92]
  wire [7:0] _tempWrData_tempMask_T_5 = reqReg_storeMask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_7 = reqReg_storeMask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_9 = reqReg_storeMask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _tempWrData_tempMask_T_11 = reqReg_storeMask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [31:0] tempWrData_tempMask = {_tempWrData_tempMask_T_11,_tempWrData_tempMask_T_9,_tempWrData_tempMask_T_7,
    _tempWrData_tempMask_T_5}; // @[Cat.scala 33:92]
  wire [31:0] _tempWrData_T = ~tempWrData_tempMask; // @[Parameters.scala 67:8]
  wire [31:0] _tempWrData_T_1 = _tempWrData_T & _GEN_35; // @[Parameters.scala 67:18]
  wire [31:0] _tempWrData_T_2 = tempWrData_tempMask & reqReg_storeData; // @[Parameters.scala 67:41]
  wire [31:0] _tempWrData_T_3 = _tempWrData_T_1 | _tempWrData_T_2; // @[Parameters.scala 67:29]
  reg [31:0] io_resp_load_bits_data_r; // @[Reg.scala 19:16]
  assign io_req_ready = state == 3'h0; // @[MSHR.scala 68:27]
  assign io_resp_load_valid = _willRespLoad_T_1 & (_T_14 | willRespLoad); // @[MSHR.scala 166:40]
  assign io_resp_load_bits_data = _T_5 ? io_tasks_refill_resp_bits_data : io_resp_load_bits_data_r; // @[MSHR.scala 167:34]
  assign io_resp_store_valid = _GEN_17 & (_T_14 | willRespStore); // @[MSHR.scala 172:40]
  assign io_tasks_refill_req_valid = _T_4 | willRefill; // @[MSHR.scala 132:52]
  assign io_tasks_refill_req_bits_addr = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[MSHR.scala 60:18]
  assign io_tasks_refill_req_bits_chosenWay = _reqReg_T ? io_req_bits_dirInfo_chosenWay : reqReg_dirInfo_chosenWay; // @[MSHR.scala 60:18]
  assign io_tasks_refill_resp_ready = 1'h1; // @[MSHR.scala 135:32]
  assign io_tasks_writeback_req_valid = _T_2 | willWriteback; // @[MSHR.scala 138:58]
  assign io_tasks_writeback_req_bits_addr = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[MSHR.scala 60:18]
  assign io_tasks_writeback_req_bits_dirtyTag = _reqReg_T ? io_req_bits_dirtyTag : reqReg_dirtyTag; // @[MSHR.scala 60:18]
  assign io_tasks_writeback_req_bits_data_0 = _reqReg_T ? io_req_bits_data_0 : reqReg_data_0; // @[MSHR.scala 60:18]
  assign io_tasks_writeback_req_bits_data_1 = _reqReg_T ? io_req_bits_data_1 : reqReg_data_1; // @[MSHR.scala 60:18]
  assign io_tasks_writeback_req_bits_data_2 = _reqReg_T ? io_req_bits_data_2 : reqReg_data_2; // @[MSHR.scala 60:18]
  assign io_tasks_writeback_req_bits_data_3 = _reqReg_T ? io_req_bits_data_3 : reqReg_data_3; // @[MSHR.scala 60:18]
  assign io_tasks_writeback_resp_ready = 1'h1; // @[MSHR.scala 142:35]
  assign io_dirWrite_req_valid = _T_9 | willWriteStore; // @[MSHR.scala 145:51]
  assign io_dirWrite_req_bits_addr = reqReg_addr; // @[MSHR.scala 146:31]
  assign io_dirWrite_req_bits_way = reqReg_dirInfo_chosenWay; // @[MSHR.scala 151:30]
  assign io_dataWrite_req_valid = _T_9 | willWriteStore; // @[MSHR.scala 154:52]
  assign io_dataWrite_req_bits_set = reqReg_addr[11:4]; // @[Parameters.scala 50:11]
  assign io_dataWrite_req_bits_data_0 = 2'h0 == _T_23 ? _tempWrData_T_3 : 32'h0; // @[MSHR.scala 159:30 160:{60,60}]
  assign io_dataWrite_req_bits_data_1 = 2'h1 == _T_23 ? _tempWrData_T_3 : 32'h0; // @[MSHR.scala 159:30 160:{60,60}]
  assign io_dataWrite_req_bits_data_2 = 2'h2 == _T_23 ? _tempWrData_T_3 : 32'h0; // @[MSHR.scala 159:30 160:{60,60}]
  assign io_dataWrite_req_bits_data_3 = 2'h3 == _T_23 ? _tempWrData_T_3 : 32'h0; // @[MSHR.scala 159:30 160:{60,60}]
  assign io_dataWrite_req_bits_blockMask = 4'h1 << reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  assign io_dataWrite_req_bits_way = reqReg_dirInfo_chosenWay; // @[MSHR.scala 157:31]
  always @(posedge clock) begin
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_addr <= io_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_dirInfo_chosenWay <= io_req_bits_dirInfo_chosenWay; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_dirtyTag <= io_req_bits_dirtyTag; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_0 <= io_req_bits_data_0; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_1 <= io_req_bits_data_1; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_2 <= io_req_bits_data_2; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_3 <= io_req_bits_data_3; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_isStore <= io_req_bits_isStore; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_storeData <= io_req_bits_storeData; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_storeMask <= io_req_bits_storeMask; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[MSHR.scala 64:24]
      state <= 3'h0; // @[MSHR.scala 64:24]
    end else if (state == 3'h4) begin // @[MSHR.scala 117:27]
      if (_T_8 | _T_13) begin // @[MSHR.scala 119:55]
        state <= 3'h0; // @[MSHR.scala 120:23]
      end else begin
        state <= 3'h4; // @[MSHR.scala 118:19]
      end
    end else if (state == 3'h3) begin // @[MSHR.scala 105:32]
      if (_T_13) begin // @[MSHR.scala 111:34]
        state <= 3'h0; // @[MSHR.scala 112:23]
      end else begin
        state <= _GEN_30;
      end
    end else if (state == 3'h2) begin // @[MSHR.scala 91:29]
      state <= _GEN_28;
    end else begin
      state <= {{1'd0}, _GEN_25};
    end
    if (_T_5) begin // @[Reg.scala 20:18]
      oldData_r <= io_tasks_refill_resp_bits_data; // @[Reg.scala 20:22]
    end
    if (_T_5) begin // @[Reg.scala 20:18]
      io_resp_load_bits_data_r <= io_tasks_refill_resp_bits_data; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reqReg_addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reqReg_dirInfo_chosenWay = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  reqReg_dirtyTag = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  reqReg_data_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reqReg_data_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reqReg_data_2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reqReg_data_3 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reqReg_isStore = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reqReg_storeData = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reqReg_storeMask = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  oldData_r = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  io_resp_load_bits_data_r = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RefillPipe_1(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [31:0]  io_req_bits_addr,
  input  [7:0]   io_req_bits_chosenWay,
  output         io_resp_valid,
  output [31:0]  io_resp_bits_data,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [127:0] io_tlbus_req_bits_size,
  output [31:0]  io_tlbus_req_bits_address,
  output         io_tlbus_resp_ready,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data,
  input          io_dirWrite_req_ready,
  output         io_dirWrite_req_valid,
  output [31:0]  io_dirWrite_req_bits_addr,
  output [7:0]   io_dirWrite_req_bits_way,
  input          io_dataWrite_req_ready,
  output         io_dataWrite_req_valid,
  output [7:0]   io_dataWrite_req_bits_set,
  output [31:0]  io_dataWrite_req_bits_data_0,
  output [31:0]  io_dataWrite_req_bits_data_1,
  output [31:0]  io_dataWrite_req_bits_data_2,
  output [31:0]  io_dataWrite_req_bits_data_3,
  output [7:0]   io_dataWrite_req_bits_way
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[RefillPipe.scala 42:24]
  wire  _io_req_ready_T = state == 2'h0; // @[RefillPipe.scala 45:27]
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] reqReg_addr; // @[Reg.scala 19:16]
  reg [7:0] reqReg_chosenWay; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  reg  reqValidReg; // @[Reg.scala 19:16]
  wire  _GEN_2 = _reqReg_T | reqValidReg; // @[Reg.scala 19:16 20:{18,22}]
  wire [3:0] dataBlockSelOH = 4'h1 << reqReg_addr[3:2]; // @[OneHot.scala 57:35]
  wire  _refillFire_T = io_tlbus_resp_ready & io_tlbus_resp_valid; // @[Decoupled.scala 51:35]
  wire  refillFire = _refillFire_T & io_tlbus_resp_bits_opcode == 3'h1; // @[RefillPipe.scala 59:41]
  wire  _T_2 = io_tlbus_req_ready & io_tlbus_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_4 = _T_2 ? 2'h2 : {{1'd0}, _reqReg_T}; // @[RefillPipe.scala 71:33 72:23]
  wire  _GEN_5 = _T_2 ? 1'h0 : _GEN_2; // @[RefillPipe.scala 71:33 73:25]
  wire [1:0] _GEN_6 = _io_req_ready_T ? _GEN_4 : 2'h0; // @[RefillPipe.scala 66:27 43:29]
  wire  _GEN_7 = _io_req_ready_T ? _GEN_5 : _GEN_2; // @[RefillPipe.scala 66:27]
  wire [1:0] _GEN_8 = _T_2 ? 2'h2 : 2'h1; // @[RefillPipe.scala 80:19 81:33 82:23]
  wire  _T_5 = state == 2'h2; // @[RefillPipe.scala 89:16]
  wire [1:0] _GEN_12 = io_resp_valid ? 2'h0 : 2'h3; // @[RefillPipe.scala 92:23 93:32 94:27]
  wire  _T_7 = state == 2'h3; // @[RefillPipe.scala 105:16]
  wire [31:0] _io_resp_bits_data_T_8 = dataBlockSelOH[0] ? io_tlbus_resp_bits_data[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_9 = dataBlockSelOH[1] ? io_tlbus_resp_bits_data[63:32] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_10 = dataBlockSelOH[2] ? io_tlbus_resp_bits_data[95:64] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_11 = dataBlockSelOH[3] ? io_tlbus_resp_bits_data[127:96] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_12 = _io_resp_bits_data_T_8 | _io_resp_bits_data_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_resp_bits_data_T_13 = _io_resp_bits_data_T_12 | _io_resp_bits_data_T_10; // @[Mux.scala 27:73]
  reg [63:0] c; // @[util.scala 162:24]
  wire [63:0] _c_T_1 = c + 64'h1; // @[util.scala 163:16]
  reg [63:0] c_1; // @[util.scala 162:24]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[util.scala 163:16]
  assign io_req_ready = state == 2'h0; // @[RefillPipe.scala 45:27]
  assign io_resp_valid = _T_7 | refillFire; // @[RefillPipe.scala 140:38]
  assign io_resp_bits_data = _io_resp_bits_data_T_13 | _io_resp_bits_data_T_11; // @[Mux.scala 27:73]
  assign io_tlbus_req_valid = _reqReg_T | reqValidReg; // @[RefillPipe.scala 50:23]
  assign io_tlbus_req_bits_size = 128'h10; // @[RefillPipe.scala 150:28]
  assign io_tlbus_req_bits_address = {_GEN_0[31:4],4'h0}; // @[Cat.scala 33:92]
  assign io_tlbus_resp_ready = io_dataWrite_req_ready & io_dirWrite_req_ready; // @[RefillPipe.scala 62:51]
  assign io_dirWrite_req_valid = refillFire & _T_5; // @[RefillPipe.scala 115:33]
  assign io_dirWrite_req_bits_addr = reqReg_addr; // @[RefillPipe.scala 117:31]
  assign io_dirWrite_req_bits_way = reqReg_chosenWay; // @[RefillPipe.scala 122:30]
  assign io_dataWrite_req_valid = refillFire & _T_5; // @[RefillPipe.scala 115:33]
  assign io_dataWrite_req_bits_set = reqReg_addr[11:4]; // @[Parameters.scala 50:11]
  assign io_dataWrite_req_bits_data_0 = io_tlbus_resp_bits_data[31:0]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_1 = io_tlbus_resp_bits_data[63:32]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_2 = io_tlbus_resp_bits_data[95:64]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_data_3 = io_tlbus_resp_bits_data[127:96]; // @[RefillPipe.scala 130:99]
  assign io_dataWrite_req_bits_way = reqReg_chosenWay; // @[RefillPipe.scala 128:31]
  always @(posedge clock) begin
    if (reset) begin // @[RefillPipe.scala 42:24]
      state <= 2'h0; // @[RefillPipe.scala 42:24]
    end else if (state == 2'h3) begin // @[RefillPipe.scala 105:27]
      state <= _GEN_12;
    end else if (state == 2'h2) begin // @[RefillPipe.scala 89:33]
      if (refillFire) begin // @[RefillPipe.scala 91:30]
        state <= _GEN_12;
      end else begin
        state <= 2'h2;
      end
    end else if (state == 2'h1) begin // @[RefillPipe.scala 79:26]
      state <= _GEN_8;
    end else begin
      state <= _GEN_6;
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_addr <= io_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_chosenWay <= io_req_bits_chosenWay; // @[Reg.scala 20:22]
    end
    if (state == 2'h1) begin // @[RefillPipe.scala 79:26]
      if (_T_2) begin // @[RefillPipe.scala 81:33]
        reqValidReg <= 1'h0; // @[RefillPipe.scala 83:25]
      end else begin
        reqValidReg <= _GEN_7;
      end
    end else begin
      reqValidReg <= _GEN_7;
    end
    if (reset) begin // @[util.scala 162:24]
      c <= 64'h0; // @[util.scala 162:24]
    end else begin
      c <= _c_T_1; // @[util.scala 163:11]
    end
    if (reset) begin // @[util.scala 162:24]
      c_1 <= 64'h0; // @[util.scala 162:24]
    end else begin
      c_1 <= _c_T_3; // @[util.scala 163:11]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [RefillPipe] req ==> addr: 0x%x size:%d\n",c,
            io_tlbus_req_bits_address,io_tlbus_req_bits_size); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (refillFire & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [RefillPipe] resp <== data: 0x%x beat: %d\n",c_1,
            io_tlbus_resp_bits_data,1'h0); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reqReg_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqReg_chosenWay = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  reqValidReg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  c = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c_1 = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLSerializer(
  input         io_in_valid,
  input  [31:0] io_in_bits_0_0,
  input  [31:0] io_in_bits_0_1,
  input  [31:0] io_in_bits_0_2,
  input  [31:0] io_in_bits_0_3,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_0,
  output [31:0] io_out_bits_1,
  output [31:0] io_out_bits_2,
  output [31:0] io_out_bits_3,
  output        io_fireAll
);
  assign io_out_valid = io_in_valid; // @[TLSerializer.scala 41:18]
  assign io_out_bits_0 = io_in_bits_0_0; // @[TLSerializer.scala 42:17]
  assign io_out_bits_1 = io_in_bits_0_1; // @[TLSerializer.scala 42:17]
  assign io_out_bits_2 = io_in_bits_0_2; // @[TLSerializer.scala 42:17]
  assign io_out_bits_3 = io_in_bits_0_3; // @[TLSerializer.scala 42:17]
  assign io_fireAll = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
endmodule
module WritebackQueue(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [31:0]  io_req_bits_addr,
  input  [19:0]  io_req_bits_dirtyTag,
  input  [31:0]  io_req_bits_data_0,
  input  [31:0]  io_req_bits_data_1,
  input  [31:0]  io_req_bits_data_2,
  input  [31:0]  io_req_bits_data_3,
  output         io_resp_valid,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [31:0]  io_tlbus_req_bits_address,
  output [127:0] io_tlbus_req_bits_data,
  output         io_tlbus_resp_ready,
  input          io_tlbus_resp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  serializer_io_in_valid; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_in_bits_0_0; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_in_bits_0_1; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_in_bits_0_2; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_in_bits_0_3; // @[WritebackQueue.scala 49:28]
  wire  serializer_io_out_ready; // @[WritebackQueue.scala 49:28]
  wire  serializer_io_out_valid; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_out_bits_0; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_out_bits_1; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_out_bits_2; // @[WritebackQueue.scala 49:28]
  wire [31:0] serializer_io_out_bits_3; // @[WritebackQueue.scala 49:28]
  wire  serializer_io_fireAll; // @[WritebackQueue.scala 49:28]
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [31:0] reqReg_addr; // @[Reg.scala 19:16]
  reg [19:0] reqReg_dirtyTag; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_0; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_1; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_2; // @[Reg.scala 19:16]
  reg [31:0] reqReg_data_3; // @[Reg.scala 19:16]
  wire [31:0] _GEN_0 = _reqReg_T ? io_req_bits_addr : reqReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire [19:0] _GEN_1 = _reqReg_T ? io_req_bits_dirtyTag : reqReg_dirtyTag; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_2 = _reqReg_T ? io_req_bits_data_0 : reqReg_data_0; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_3 = _reqReg_T ? io_req_bits_data_1 : reqReg_data_1; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_4 = _reqReg_T ? io_req_bits_data_2 : reqReg_data_2; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_5 = _reqReg_T ? io_req_bits_data_3 : reqReg_data_3; // @[Reg.scala 19:16 20:{18,22}]
  wire [19:0] req_dirtyTag = _reqReg_T ? io_req_bits_dirtyTag : reqReg_dirtyTag; // @[WritebackQueue.scala 43:18]
  reg  reqValidReg; // @[Reg.scala 19:16]
  wire  _GEN_6 = _reqReg_T | reqValidReg; // @[Reg.scala 19:16 20:{18,22}]
  wire [127:0] _T = {_GEN_5,_GEN_4,_GEN_3,_GEN_2}; // @[WritebackQueue.scala 51:47]
  reg [1:0] state; // @[WritebackQueue.scala 53:24]
  wire  _io_req_ready_T = state == 2'h0; // @[WritebackQueue.scala 56:27]
  wire  _GEN_8 = _io_req_ready_T & _reqReg_T; // @[WritebackQueue.scala 58:27 54:29]
  wire [1:0] _GEN_9 = serializer_io_fireAll ? 2'h2 : 2'h1; // @[WritebackQueue.scala 66:19 67:37 68:23]
  wire  _GEN_10 = serializer_io_fireAll ? 1'h0 : _GEN_6; // @[WritebackQueue.scala 67:37 70:25]
  wire  _GEN_12 = state == 2'h1 ? _GEN_10 : _GEN_6; // @[WritebackQueue.scala 65:34]
  wire  _T_8 = state == 2'h2; // @[WritebackQueue.scala 74:16]
  wire  _T_9 = io_tlbus_resp_ready & io_tlbus_resp_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_13 = io_resp_valid ? 2'h0 : 2'h3; // @[WritebackQueue.scala 77:23 79:32 80:27]
  wire  _T_11 = state == 2'h3; // @[WritebackQueue.scala 85:16]
  wire [63:0] io_tlbus_req_bits_data_lo = {serializer_io_out_bits_1,serializer_io_out_bits_0}; // @[WritebackQueue.scala 103:54]
  wire [63:0] io_tlbus_req_bits_data_hi = {serializer_io_out_bits_3,serializer_io_out_bits_2}; // @[WritebackQueue.scala 103:54]
  wire [7:0] dirtySet = _GEN_0[11:4]; // @[Parameters.scala 50:11]
  wire [31:0] writebackAddr = {_GEN_1,dirtySet,4'h0}; // @[Cat.scala 33:92]
  wire [32:0] _io_tlbus_req_bits_address_T_1 = {{1'd0}, writebackAddr}; // @[WritebackQueue.scala 110:49]
  TLSerializer serializer ( // @[WritebackQueue.scala 49:28]
    .io_in_valid(serializer_io_in_valid),
    .io_in_bits_0_0(serializer_io_in_bits_0_0),
    .io_in_bits_0_1(serializer_io_in_bits_0_1),
    .io_in_bits_0_2(serializer_io_in_bits_0_2),
    .io_in_bits_0_3(serializer_io_in_bits_0_3),
    .io_out_ready(serializer_io_out_ready),
    .io_out_valid(serializer_io_out_valid),
    .io_out_bits_0(serializer_io_out_bits_0),
    .io_out_bits_1(serializer_io_out_bits_1),
    .io_out_bits_2(serializer_io_out_bits_2),
    .io_out_bits_3(serializer_io_out_bits_3),
    .io_fireAll(serializer_io_fireAll)
  );
  assign io_req_ready = state == 2'h0; // @[WritebackQueue.scala 56:27]
  assign io_resp_valid = _T_11 | _T_9 & _T_8; // @[WritebackQueue.scala 96:38]
  assign io_tlbus_req_valid = serializer_io_out_valid; // @[WritebackQueue.scala 101:24]
  assign io_tlbus_req_bits_address = _io_tlbus_req_bits_address_T_1[31:0]; // @[WritebackQueue.scala 110:49]
  assign io_tlbus_req_bits_data = {io_tlbus_req_bits_data_hi,io_tlbus_req_bits_data_lo}; // @[WritebackQueue.scala 103:54]
  assign io_tlbus_resp_ready = 1'h1; // @[WritebackQueue.scala 98:25]
  assign serializer_io_in_valid = _reqReg_T | reqValidReg; // @[WritebackQueue.scala 45:23]
  assign serializer_io_in_bits_0_0 = _T[31:0]; // @[WritebackQueue.scala 51:47]
  assign serializer_io_in_bits_0_1 = _T[63:32]; // @[WritebackQueue.scala 51:47]
  assign serializer_io_in_bits_0_2 = _T[95:64]; // @[WritebackQueue.scala 51:47]
  assign serializer_io_in_bits_0_3 = _T[127:96]; // @[WritebackQueue.scala 51:47]
  assign serializer_io_out_ready = io_tlbus_req_ready; // @[WritebackQueue.scala 100:29]
  always @(posedge clock) begin
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_addr <= io_req_bits_addr; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_dirtyTag <= io_req_bits_dirtyTag; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_0 <= io_req_bits_data_0; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_1 <= io_req_bits_data_1; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_2 <= io_req_bits_data_2; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data_3 <= io_req_bits_data_3; // @[Reg.scala 20:22]
    end
    if (state == 2'h3) begin // @[WritebackQueue.scala 85:27]
      if (io_resp_valid) begin // @[WritebackQueue.scala 87:28]
        reqValidReg <= 1'h0; // @[WritebackQueue.scala 90:25]
      end else begin
        reqValidReg <= _GEN_12;
      end
    end else begin
      reqValidReg <= _GEN_12;
    end
    if (reset) begin // @[WritebackQueue.scala 53:24]
      state <= 2'h0; // @[WritebackQueue.scala 53:24]
    end else if (state == 2'h3) begin // @[WritebackQueue.scala 85:27]
      state <= _GEN_13;
    end else if (state == 2'h2) begin // @[WritebackQueue.scala 74:32]
      if (_T_9) begin // @[WritebackQueue.scala 76:34]
        state <= _GEN_13;
      end else begin
        state <= 2'h2; // @[WritebackQueue.scala 75:19]
      end
    end else if (state == 2'h1) begin // @[WritebackQueue.scala 65:34]
      state <= _GEN_9;
    end else begin
      state <= {{1'd0}, _GEN_8};
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reqReg_addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reqReg_dirtyTag = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  reqReg_data_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reqReg_data_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reqReg_data_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reqReg_data_3 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reqValidReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BankRAM_2P_80(
  input         clock,
  input         reset,
  input  [7:0]  io_r_addr,
  output [31:0] io_r_data,
  input         io_w_en,
  input  [7:0]  io_w_addr,
  input  [31:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:255]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_129_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_130_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_131_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_132_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_133_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_134_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_135_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_136_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_137_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_138_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_139_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_140_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_141_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_142_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_143_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_144_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_145_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_146_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_147_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_148_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_149_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_150_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_151_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_152_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_153_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_154_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_155_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_156_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_157_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_158_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_159_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_160_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_161_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_162_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_163_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_164_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_165_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_166_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_167_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_168_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_169_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_170_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_171_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_172_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_173_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_174_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_175_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_176_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_177_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_178_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_179_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_180_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_181_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_182_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_183_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_184_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_185_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_186_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_187_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_188_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_189_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_190_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_191_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_192_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_193_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_194_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_195_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_196_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_197_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_198_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_199_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_200_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_201_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_202_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_203_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_204_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_205_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_206_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_207_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_208_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_209_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_210_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_211_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_212_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_213_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_214_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_215_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_216_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_217_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_218_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_219_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_220_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_221_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_222_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_223_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_224_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_225_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_226_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_227_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_228_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_229_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_230_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_231_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_232_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_233_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_234_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_235_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_236_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_237_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_238_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_239_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_240_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_241_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_242_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_243_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_244_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_245_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_246_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_247_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_248_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_249_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_250_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_251_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_252_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_253_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_254_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_255_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_en; // @[SRAM_1.scala 63:26]
  wire [31:0] mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_256_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [7:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 32'h0;
  assign mem_MPORT_addr = 8'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 32'h0;
  assign mem_MPORT_1_addr = 8'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 32'h0;
  assign mem_MPORT_2_addr = 8'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 32'h0;
  assign mem_MPORT_3_addr = 8'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 32'h0;
  assign mem_MPORT_4_addr = 8'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 32'h0;
  assign mem_MPORT_5_addr = 8'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 32'h0;
  assign mem_MPORT_6_addr = 8'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 32'h0;
  assign mem_MPORT_7_addr = 8'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 32'h0;
  assign mem_MPORT_8_addr = 8'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 32'h0;
  assign mem_MPORT_9_addr = 8'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 32'h0;
  assign mem_MPORT_10_addr = 8'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 32'h0;
  assign mem_MPORT_11_addr = 8'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 32'h0;
  assign mem_MPORT_12_addr = 8'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 32'h0;
  assign mem_MPORT_13_addr = 8'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 32'h0;
  assign mem_MPORT_14_addr = 8'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 32'h0;
  assign mem_MPORT_15_addr = 8'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 32'h0;
  assign mem_MPORT_16_addr = 8'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 32'h0;
  assign mem_MPORT_17_addr = 8'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 32'h0;
  assign mem_MPORT_18_addr = 8'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 32'h0;
  assign mem_MPORT_19_addr = 8'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 32'h0;
  assign mem_MPORT_20_addr = 8'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 32'h0;
  assign mem_MPORT_21_addr = 8'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 32'h0;
  assign mem_MPORT_22_addr = 8'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 32'h0;
  assign mem_MPORT_23_addr = 8'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 32'h0;
  assign mem_MPORT_24_addr = 8'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 32'h0;
  assign mem_MPORT_25_addr = 8'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 32'h0;
  assign mem_MPORT_26_addr = 8'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 32'h0;
  assign mem_MPORT_27_addr = 8'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 32'h0;
  assign mem_MPORT_28_addr = 8'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 32'h0;
  assign mem_MPORT_29_addr = 8'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 32'h0;
  assign mem_MPORT_30_addr = 8'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 32'h0;
  assign mem_MPORT_31_addr = 8'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 32'h0;
  assign mem_MPORT_32_addr = 8'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 32'h0;
  assign mem_MPORT_33_addr = 8'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 32'h0;
  assign mem_MPORT_34_addr = 8'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 32'h0;
  assign mem_MPORT_35_addr = 8'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 32'h0;
  assign mem_MPORT_36_addr = 8'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 32'h0;
  assign mem_MPORT_37_addr = 8'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 32'h0;
  assign mem_MPORT_38_addr = 8'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 32'h0;
  assign mem_MPORT_39_addr = 8'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 32'h0;
  assign mem_MPORT_40_addr = 8'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 32'h0;
  assign mem_MPORT_41_addr = 8'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 32'h0;
  assign mem_MPORT_42_addr = 8'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 32'h0;
  assign mem_MPORT_43_addr = 8'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 32'h0;
  assign mem_MPORT_44_addr = 8'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 32'h0;
  assign mem_MPORT_45_addr = 8'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 32'h0;
  assign mem_MPORT_46_addr = 8'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 32'h0;
  assign mem_MPORT_47_addr = 8'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 32'h0;
  assign mem_MPORT_48_addr = 8'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 32'h0;
  assign mem_MPORT_49_addr = 8'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 32'h0;
  assign mem_MPORT_50_addr = 8'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 32'h0;
  assign mem_MPORT_51_addr = 8'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 32'h0;
  assign mem_MPORT_52_addr = 8'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 32'h0;
  assign mem_MPORT_53_addr = 8'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 32'h0;
  assign mem_MPORT_54_addr = 8'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 32'h0;
  assign mem_MPORT_55_addr = 8'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 32'h0;
  assign mem_MPORT_56_addr = 8'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 32'h0;
  assign mem_MPORT_57_addr = 8'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 32'h0;
  assign mem_MPORT_58_addr = 8'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 32'h0;
  assign mem_MPORT_59_addr = 8'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 32'h0;
  assign mem_MPORT_60_addr = 8'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 32'h0;
  assign mem_MPORT_61_addr = 8'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 32'h0;
  assign mem_MPORT_62_addr = 8'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 32'h0;
  assign mem_MPORT_63_addr = 8'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 32'h0;
  assign mem_MPORT_64_addr = 8'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 32'h0;
  assign mem_MPORT_65_addr = 8'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 32'h0;
  assign mem_MPORT_66_addr = 8'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 32'h0;
  assign mem_MPORT_67_addr = 8'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 32'h0;
  assign mem_MPORT_68_addr = 8'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 32'h0;
  assign mem_MPORT_69_addr = 8'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 32'h0;
  assign mem_MPORT_70_addr = 8'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 32'h0;
  assign mem_MPORT_71_addr = 8'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 32'h0;
  assign mem_MPORT_72_addr = 8'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 32'h0;
  assign mem_MPORT_73_addr = 8'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 32'h0;
  assign mem_MPORT_74_addr = 8'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 32'h0;
  assign mem_MPORT_75_addr = 8'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 32'h0;
  assign mem_MPORT_76_addr = 8'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 32'h0;
  assign mem_MPORT_77_addr = 8'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 32'h0;
  assign mem_MPORT_78_addr = 8'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 32'h0;
  assign mem_MPORT_79_addr = 8'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 32'h0;
  assign mem_MPORT_80_addr = 8'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 32'h0;
  assign mem_MPORT_81_addr = 8'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 32'h0;
  assign mem_MPORT_82_addr = 8'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 32'h0;
  assign mem_MPORT_83_addr = 8'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 32'h0;
  assign mem_MPORT_84_addr = 8'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 32'h0;
  assign mem_MPORT_85_addr = 8'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 32'h0;
  assign mem_MPORT_86_addr = 8'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 32'h0;
  assign mem_MPORT_87_addr = 8'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 32'h0;
  assign mem_MPORT_88_addr = 8'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 32'h0;
  assign mem_MPORT_89_addr = 8'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 32'h0;
  assign mem_MPORT_90_addr = 8'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 32'h0;
  assign mem_MPORT_91_addr = 8'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 32'h0;
  assign mem_MPORT_92_addr = 8'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 32'h0;
  assign mem_MPORT_93_addr = 8'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 32'h0;
  assign mem_MPORT_94_addr = 8'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 32'h0;
  assign mem_MPORT_95_addr = 8'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 32'h0;
  assign mem_MPORT_96_addr = 8'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 32'h0;
  assign mem_MPORT_97_addr = 8'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 32'h0;
  assign mem_MPORT_98_addr = 8'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 32'h0;
  assign mem_MPORT_99_addr = 8'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 32'h0;
  assign mem_MPORT_100_addr = 8'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 32'h0;
  assign mem_MPORT_101_addr = 8'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 32'h0;
  assign mem_MPORT_102_addr = 8'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 32'h0;
  assign mem_MPORT_103_addr = 8'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 32'h0;
  assign mem_MPORT_104_addr = 8'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 32'h0;
  assign mem_MPORT_105_addr = 8'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 32'h0;
  assign mem_MPORT_106_addr = 8'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 32'h0;
  assign mem_MPORT_107_addr = 8'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 32'h0;
  assign mem_MPORT_108_addr = 8'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 32'h0;
  assign mem_MPORT_109_addr = 8'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 32'h0;
  assign mem_MPORT_110_addr = 8'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 32'h0;
  assign mem_MPORT_111_addr = 8'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 32'h0;
  assign mem_MPORT_112_addr = 8'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 32'h0;
  assign mem_MPORT_113_addr = 8'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 32'h0;
  assign mem_MPORT_114_addr = 8'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 32'h0;
  assign mem_MPORT_115_addr = 8'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 32'h0;
  assign mem_MPORT_116_addr = 8'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 32'h0;
  assign mem_MPORT_117_addr = 8'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 32'h0;
  assign mem_MPORT_118_addr = 8'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 32'h0;
  assign mem_MPORT_119_addr = 8'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 32'h0;
  assign mem_MPORT_120_addr = 8'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 32'h0;
  assign mem_MPORT_121_addr = 8'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 32'h0;
  assign mem_MPORT_122_addr = 8'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 32'h0;
  assign mem_MPORT_123_addr = 8'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 32'h0;
  assign mem_MPORT_124_addr = 8'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 32'h0;
  assign mem_MPORT_125_addr = 8'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 32'h0;
  assign mem_MPORT_126_addr = 8'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 32'h0;
  assign mem_MPORT_127_addr = 8'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 32'h0;
  assign mem_MPORT_128_addr = 8'h80;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = reset;
  assign mem_MPORT_129_data = 32'h0;
  assign mem_MPORT_129_addr = 8'h81;
  assign mem_MPORT_129_mask = 1'h1;
  assign mem_MPORT_129_en = reset;
  assign mem_MPORT_130_data = 32'h0;
  assign mem_MPORT_130_addr = 8'h82;
  assign mem_MPORT_130_mask = 1'h1;
  assign mem_MPORT_130_en = reset;
  assign mem_MPORT_131_data = 32'h0;
  assign mem_MPORT_131_addr = 8'h83;
  assign mem_MPORT_131_mask = 1'h1;
  assign mem_MPORT_131_en = reset;
  assign mem_MPORT_132_data = 32'h0;
  assign mem_MPORT_132_addr = 8'h84;
  assign mem_MPORT_132_mask = 1'h1;
  assign mem_MPORT_132_en = reset;
  assign mem_MPORT_133_data = 32'h0;
  assign mem_MPORT_133_addr = 8'h85;
  assign mem_MPORT_133_mask = 1'h1;
  assign mem_MPORT_133_en = reset;
  assign mem_MPORT_134_data = 32'h0;
  assign mem_MPORT_134_addr = 8'h86;
  assign mem_MPORT_134_mask = 1'h1;
  assign mem_MPORT_134_en = reset;
  assign mem_MPORT_135_data = 32'h0;
  assign mem_MPORT_135_addr = 8'h87;
  assign mem_MPORT_135_mask = 1'h1;
  assign mem_MPORT_135_en = reset;
  assign mem_MPORT_136_data = 32'h0;
  assign mem_MPORT_136_addr = 8'h88;
  assign mem_MPORT_136_mask = 1'h1;
  assign mem_MPORT_136_en = reset;
  assign mem_MPORT_137_data = 32'h0;
  assign mem_MPORT_137_addr = 8'h89;
  assign mem_MPORT_137_mask = 1'h1;
  assign mem_MPORT_137_en = reset;
  assign mem_MPORT_138_data = 32'h0;
  assign mem_MPORT_138_addr = 8'h8a;
  assign mem_MPORT_138_mask = 1'h1;
  assign mem_MPORT_138_en = reset;
  assign mem_MPORT_139_data = 32'h0;
  assign mem_MPORT_139_addr = 8'h8b;
  assign mem_MPORT_139_mask = 1'h1;
  assign mem_MPORT_139_en = reset;
  assign mem_MPORT_140_data = 32'h0;
  assign mem_MPORT_140_addr = 8'h8c;
  assign mem_MPORT_140_mask = 1'h1;
  assign mem_MPORT_140_en = reset;
  assign mem_MPORT_141_data = 32'h0;
  assign mem_MPORT_141_addr = 8'h8d;
  assign mem_MPORT_141_mask = 1'h1;
  assign mem_MPORT_141_en = reset;
  assign mem_MPORT_142_data = 32'h0;
  assign mem_MPORT_142_addr = 8'h8e;
  assign mem_MPORT_142_mask = 1'h1;
  assign mem_MPORT_142_en = reset;
  assign mem_MPORT_143_data = 32'h0;
  assign mem_MPORT_143_addr = 8'h8f;
  assign mem_MPORT_143_mask = 1'h1;
  assign mem_MPORT_143_en = reset;
  assign mem_MPORT_144_data = 32'h0;
  assign mem_MPORT_144_addr = 8'h90;
  assign mem_MPORT_144_mask = 1'h1;
  assign mem_MPORT_144_en = reset;
  assign mem_MPORT_145_data = 32'h0;
  assign mem_MPORT_145_addr = 8'h91;
  assign mem_MPORT_145_mask = 1'h1;
  assign mem_MPORT_145_en = reset;
  assign mem_MPORT_146_data = 32'h0;
  assign mem_MPORT_146_addr = 8'h92;
  assign mem_MPORT_146_mask = 1'h1;
  assign mem_MPORT_146_en = reset;
  assign mem_MPORT_147_data = 32'h0;
  assign mem_MPORT_147_addr = 8'h93;
  assign mem_MPORT_147_mask = 1'h1;
  assign mem_MPORT_147_en = reset;
  assign mem_MPORT_148_data = 32'h0;
  assign mem_MPORT_148_addr = 8'h94;
  assign mem_MPORT_148_mask = 1'h1;
  assign mem_MPORT_148_en = reset;
  assign mem_MPORT_149_data = 32'h0;
  assign mem_MPORT_149_addr = 8'h95;
  assign mem_MPORT_149_mask = 1'h1;
  assign mem_MPORT_149_en = reset;
  assign mem_MPORT_150_data = 32'h0;
  assign mem_MPORT_150_addr = 8'h96;
  assign mem_MPORT_150_mask = 1'h1;
  assign mem_MPORT_150_en = reset;
  assign mem_MPORT_151_data = 32'h0;
  assign mem_MPORT_151_addr = 8'h97;
  assign mem_MPORT_151_mask = 1'h1;
  assign mem_MPORT_151_en = reset;
  assign mem_MPORT_152_data = 32'h0;
  assign mem_MPORT_152_addr = 8'h98;
  assign mem_MPORT_152_mask = 1'h1;
  assign mem_MPORT_152_en = reset;
  assign mem_MPORT_153_data = 32'h0;
  assign mem_MPORT_153_addr = 8'h99;
  assign mem_MPORT_153_mask = 1'h1;
  assign mem_MPORT_153_en = reset;
  assign mem_MPORT_154_data = 32'h0;
  assign mem_MPORT_154_addr = 8'h9a;
  assign mem_MPORT_154_mask = 1'h1;
  assign mem_MPORT_154_en = reset;
  assign mem_MPORT_155_data = 32'h0;
  assign mem_MPORT_155_addr = 8'h9b;
  assign mem_MPORT_155_mask = 1'h1;
  assign mem_MPORT_155_en = reset;
  assign mem_MPORT_156_data = 32'h0;
  assign mem_MPORT_156_addr = 8'h9c;
  assign mem_MPORT_156_mask = 1'h1;
  assign mem_MPORT_156_en = reset;
  assign mem_MPORT_157_data = 32'h0;
  assign mem_MPORT_157_addr = 8'h9d;
  assign mem_MPORT_157_mask = 1'h1;
  assign mem_MPORT_157_en = reset;
  assign mem_MPORT_158_data = 32'h0;
  assign mem_MPORT_158_addr = 8'h9e;
  assign mem_MPORT_158_mask = 1'h1;
  assign mem_MPORT_158_en = reset;
  assign mem_MPORT_159_data = 32'h0;
  assign mem_MPORT_159_addr = 8'h9f;
  assign mem_MPORT_159_mask = 1'h1;
  assign mem_MPORT_159_en = reset;
  assign mem_MPORT_160_data = 32'h0;
  assign mem_MPORT_160_addr = 8'ha0;
  assign mem_MPORT_160_mask = 1'h1;
  assign mem_MPORT_160_en = reset;
  assign mem_MPORT_161_data = 32'h0;
  assign mem_MPORT_161_addr = 8'ha1;
  assign mem_MPORT_161_mask = 1'h1;
  assign mem_MPORT_161_en = reset;
  assign mem_MPORT_162_data = 32'h0;
  assign mem_MPORT_162_addr = 8'ha2;
  assign mem_MPORT_162_mask = 1'h1;
  assign mem_MPORT_162_en = reset;
  assign mem_MPORT_163_data = 32'h0;
  assign mem_MPORT_163_addr = 8'ha3;
  assign mem_MPORT_163_mask = 1'h1;
  assign mem_MPORT_163_en = reset;
  assign mem_MPORT_164_data = 32'h0;
  assign mem_MPORT_164_addr = 8'ha4;
  assign mem_MPORT_164_mask = 1'h1;
  assign mem_MPORT_164_en = reset;
  assign mem_MPORT_165_data = 32'h0;
  assign mem_MPORT_165_addr = 8'ha5;
  assign mem_MPORT_165_mask = 1'h1;
  assign mem_MPORT_165_en = reset;
  assign mem_MPORT_166_data = 32'h0;
  assign mem_MPORT_166_addr = 8'ha6;
  assign mem_MPORT_166_mask = 1'h1;
  assign mem_MPORT_166_en = reset;
  assign mem_MPORT_167_data = 32'h0;
  assign mem_MPORT_167_addr = 8'ha7;
  assign mem_MPORT_167_mask = 1'h1;
  assign mem_MPORT_167_en = reset;
  assign mem_MPORT_168_data = 32'h0;
  assign mem_MPORT_168_addr = 8'ha8;
  assign mem_MPORT_168_mask = 1'h1;
  assign mem_MPORT_168_en = reset;
  assign mem_MPORT_169_data = 32'h0;
  assign mem_MPORT_169_addr = 8'ha9;
  assign mem_MPORT_169_mask = 1'h1;
  assign mem_MPORT_169_en = reset;
  assign mem_MPORT_170_data = 32'h0;
  assign mem_MPORT_170_addr = 8'haa;
  assign mem_MPORT_170_mask = 1'h1;
  assign mem_MPORT_170_en = reset;
  assign mem_MPORT_171_data = 32'h0;
  assign mem_MPORT_171_addr = 8'hab;
  assign mem_MPORT_171_mask = 1'h1;
  assign mem_MPORT_171_en = reset;
  assign mem_MPORT_172_data = 32'h0;
  assign mem_MPORT_172_addr = 8'hac;
  assign mem_MPORT_172_mask = 1'h1;
  assign mem_MPORT_172_en = reset;
  assign mem_MPORT_173_data = 32'h0;
  assign mem_MPORT_173_addr = 8'had;
  assign mem_MPORT_173_mask = 1'h1;
  assign mem_MPORT_173_en = reset;
  assign mem_MPORT_174_data = 32'h0;
  assign mem_MPORT_174_addr = 8'hae;
  assign mem_MPORT_174_mask = 1'h1;
  assign mem_MPORT_174_en = reset;
  assign mem_MPORT_175_data = 32'h0;
  assign mem_MPORT_175_addr = 8'haf;
  assign mem_MPORT_175_mask = 1'h1;
  assign mem_MPORT_175_en = reset;
  assign mem_MPORT_176_data = 32'h0;
  assign mem_MPORT_176_addr = 8'hb0;
  assign mem_MPORT_176_mask = 1'h1;
  assign mem_MPORT_176_en = reset;
  assign mem_MPORT_177_data = 32'h0;
  assign mem_MPORT_177_addr = 8'hb1;
  assign mem_MPORT_177_mask = 1'h1;
  assign mem_MPORT_177_en = reset;
  assign mem_MPORT_178_data = 32'h0;
  assign mem_MPORT_178_addr = 8'hb2;
  assign mem_MPORT_178_mask = 1'h1;
  assign mem_MPORT_178_en = reset;
  assign mem_MPORT_179_data = 32'h0;
  assign mem_MPORT_179_addr = 8'hb3;
  assign mem_MPORT_179_mask = 1'h1;
  assign mem_MPORT_179_en = reset;
  assign mem_MPORT_180_data = 32'h0;
  assign mem_MPORT_180_addr = 8'hb4;
  assign mem_MPORT_180_mask = 1'h1;
  assign mem_MPORT_180_en = reset;
  assign mem_MPORT_181_data = 32'h0;
  assign mem_MPORT_181_addr = 8'hb5;
  assign mem_MPORT_181_mask = 1'h1;
  assign mem_MPORT_181_en = reset;
  assign mem_MPORT_182_data = 32'h0;
  assign mem_MPORT_182_addr = 8'hb6;
  assign mem_MPORT_182_mask = 1'h1;
  assign mem_MPORT_182_en = reset;
  assign mem_MPORT_183_data = 32'h0;
  assign mem_MPORT_183_addr = 8'hb7;
  assign mem_MPORT_183_mask = 1'h1;
  assign mem_MPORT_183_en = reset;
  assign mem_MPORT_184_data = 32'h0;
  assign mem_MPORT_184_addr = 8'hb8;
  assign mem_MPORT_184_mask = 1'h1;
  assign mem_MPORT_184_en = reset;
  assign mem_MPORT_185_data = 32'h0;
  assign mem_MPORT_185_addr = 8'hb9;
  assign mem_MPORT_185_mask = 1'h1;
  assign mem_MPORT_185_en = reset;
  assign mem_MPORT_186_data = 32'h0;
  assign mem_MPORT_186_addr = 8'hba;
  assign mem_MPORT_186_mask = 1'h1;
  assign mem_MPORT_186_en = reset;
  assign mem_MPORT_187_data = 32'h0;
  assign mem_MPORT_187_addr = 8'hbb;
  assign mem_MPORT_187_mask = 1'h1;
  assign mem_MPORT_187_en = reset;
  assign mem_MPORT_188_data = 32'h0;
  assign mem_MPORT_188_addr = 8'hbc;
  assign mem_MPORT_188_mask = 1'h1;
  assign mem_MPORT_188_en = reset;
  assign mem_MPORT_189_data = 32'h0;
  assign mem_MPORT_189_addr = 8'hbd;
  assign mem_MPORT_189_mask = 1'h1;
  assign mem_MPORT_189_en = reset;
  assign mem_MPORT_190_data = 32'h0;
  assign mem_MPORT_190_addr = 8'hbe;
  assign mem_MPORT_190_mask = 1'h1;
  assign mem_MPORT_190_en = reset;
  assign mem_MPORT_191_data = 32'h0;
  assign mem_MPORT_191_addr = 8'hbf;
  assign mem_MPORT_191_mask = 1'h1;
  assign mem_MPORT_191_en = reset;
  assign mem_MPORT_192_data = 32'h0;
  assign mem_MPORT_192_addr = 8'hc0;
  assign mem_MPORT_192_mask = 1'h1;
  assign mem_MPORT_192_en = reset;
  assign mem_MPORT_193_data = 32'h0;
  assign mem_MPORT_193_addr = 8'hc1;
  assign mem_MPORT_193_mask = 1'h1;
  assign mem_MPORT_193_en = reset;
  assign mem_MPORT_194_data = 32'h0;
  assign mem_MPORT_194_addr = 8'hc2;
  assign mem_MPORT_194_mask = 1'h1;
  assign mem_MPORT_194_en = reset;
  assign mem_MPORT_195_data = 32'h0;
  assign mem_MPORT_195_addr = 8'hc3;
  assign mem_MPORT_195_mask = 1'h1;
  assign mem_MPORT_195_en = reset;
  assign mem_MPORT_196_data = 32'h0;
  assign mem_MPORT_196_addr = 8'hc4;
  assign mem_MPORT_196_mask = 1'h1;
  assign mem_MPORT_196_en = reset;
  assign mem_MPORT_197_data = 32'h0;
  assign mem_MPORT_197_addr = 8'hc5;
  assign mem_MPORT_197_mask = 1'h1;
  assign mem_MPORT_197_en = reset;
  assign mem_MPORT_198_data = 32'h0;
  assign mem_MPORT_198_addr = 8'hc6;
  assign mem_MPORT_198_mask = 1'h1;
  assign mem_MPORT_198_en = reset;
  assign mem_MPORT_199_data = 32'h0;
  assign mem_MPORT_199_addr = 8'hc7;
  assign mem_MPORT_199_mask = 1'h1;
  assign mem_MPORT_199_en = reset;
  assign mem_MPORT_200_data = 32'h0;
  assign mem_MPORT_200_addr = 8'hc8;
  assign mem_MPORT_200_mask = 1'h1;
  assign mem_MPORT_200_en = reset;
  assign mem_MPORT_201_data = 32'h0;
  assign mem_MPORT_201_addr = 8'hc9;
  assign mem_MPORT_201_mask = 1'h1;
  assign mem_MPORT_201_en = reset;
  assign mem_MPORT_202_data = 32'h0;
  assign mem_MPORT_202_addr = 8'hca;
  assign mem_MPORT_202_mask = 1'h1;
  assign mem_MPORT_202_en = reset;
  assign mem_MPORT_203_data = 32'h0;
  assign mem_MPORT_203_addr = 8'hcb;
  assign mem_MPORT_203_mask = 1'h1;
  assign mem_MPORT_203_en = reset;
  assign mem_MPORT_204_data = 32'h0;
  assign mem_MPORT_204_addr = 8'hcc;
  assign mem_MPORT_204_mask = 1'h1;
  assign mem_MPORT_204_en = reset;
  assign mem_MPORT_205_data = 32'h0;
  assign mem_MPORT_205_addr = 8'hcd;
  assign mem_MPORT_205_mask = 1'h1;
  assign mem_MPORT_205_en = reset;
  assign mem_MPORT_206_data = 32'h0;
  assign mem_MPORT_206_addr = 8'hce;
  assign mem_MPORT_206_mask = 1'h1;
  assign mem_MPORT_206_en = reset;
  assign mem_MPORT_207_data = 32'h0;
  assign mem_MPORT_207_addr = 8'hcf;
  assign mem_MPORT_207_mask = 1'h1;
  assign mem_MPORT_207_en = reset;
  assign mem_MPORT_208_data = 32'h0;
  assign mem_MPORT_208_addr = 8'hd0;
  assign mem_MPORT_208_mask = 1'h1;
  assign mem_MPORT_208_en = reset;
  assign mem_MPORT_209_data = 32'h0;
  assign mem_MPORT_209_addr = 8'hd1;
  assign mem_MPORT_209_mask = 1'h1;
  assign mem_MPORT_209_en = reset;
  assign mem_MPORT_210_data = 32'h0;
  assign mem_MPORT_210_addr = 8'hd2;
  assign mem_MPORT_210_mask = 1'h1;
  assign mem_MPORT_210_en = reset;
  assign mem_MPORT_211_data = 32'h0;
  assign mem_MPORT_211_addr = 8'hd3;
  assign mem_MPORT_211_mask = 1'h1;
  assign mem_MPORT_211_en = reset;
  assign mem_MPORT_212_data = 32'h0;
  assign mem_MPORT_212_addr = 8'hd4;
  assign mem_MPORT_212_mask = 1'h1;
  assign mem_MPORT_212_en = reset;
  assign mem_MPORT_213_data = 32'h0;
  assign mem_MPORT_213_addr = 8'hd5;
  assign mem_MPORT_213_mask = 1'h1;
  assign mem_MPORT_213_en = reset;
  assign mem_MPORT_214_data = 32'h0;
  assign mem_MPORT_214_addr = 8'hd6;
  assign mem_MPORT_214_mask = 1'h1;
  assign mem_MPORT_214_en = reset;
  assign mem_MPORT_215_data = 32'h0;
  assign mem_MPORT_215_addr = 8'hd7;
  assign mem_MPORT_215_mask = 1'h1;
  assign mem_MPORT_215_en = reset;
  assign mem_MPORT_216_data = 32'h0;
  assign mem_MPORT_216_addr = 8'hd8;
  assign mem_MPORT_216_mask = 1'h1;
  assign mem_MPORT_216_en = reset;
  assign mem_MPORT_217_data = 32'h0;
  assign mem_MPORT_217_addr = 8'hd9;
  assign mem_MPORT_217_mask = 1'h1;
  assign mem_MPORT_217_en = reset;
  assign mem_MPORT_218_data = 32'h0;
  assign mem_MPORT_218_addr = 8'hda;
  assign mem_MPORT_218_mask = 1'h1;
  assign mem_MPORT_218_en = reset;
  assign mem_MPORT_219_data = 32'h0;
  assign mem_MPORT_219_addr = 8'hdb;
  assign mem_MPORT_219_mask = 1'h1;
  assign mem_MPORT_219_en = reset;
  assign mem_MPORT_220_data = 32'h0;
  assign mem_MPORT_220_addr = 8'hdc;
  assign mem_MPORT_220_mask = 1'h1;
  assign mem_MPORT_220_en = reset;
  assign mem_MPORT_221_data = 32'h0;
  assign mem_MPORT_221_addr = 8'hdd;
  assign mem_MPORT_221_mask = 1'h1;
  assign mem_MPORT_221_en = reset;
  assign mem_MPORT_222_data = 32'h0;
  assign mem_MPORT_222_addr = 8'hde;
  assign mem_MPORT_222_mask = 1'h1;
  assign mem_MPORT_222_en = reset;
  assign mem_MPORT_223_data = 32'h0;
  assign mem_MPORT_223_addr = 8'hdf;
  assign mem_MPORT_223_mask = 1'h1;
  assign mem_MPORT_223_en = reset;
  assign mem_MPORT_224_data = 32'h0;
  assign mem_MPORT_224_addr = 8'he0;
  assign mem_MPORT_224_mask = 1'h1;
  assign mem_MPORT_224_en = reset;
  assign mem_MPORT_225_data = 32'h0;
  assign mem_MPORT_225_addr = 8'he1;
  assign mem_MPORT_225_mask = 1'h1;
  assign mem_MPORT_225_en = reset;
  assign mem_MPORT_226_data = 32'h0;
  assign mem_MPORT_226_addr = 8'he2;
  assign mem_MPORT_226_mask = 1'h1;
  assign mem_MPORT_226_en = reset;
  assign mem_MPORT_227_data = 32'h0;
  assign mem_MPORT_227_addr = 8'he3;
  assign mem_MPORT_227_mask = 1'h1;
  assign mem_MPORT_227_en = reset;
  assign mem_MPORT_228_data = 32'h0;
  assign mem_MPORT_228_addr = 8'he4;
  assign mem_MPORT_228_mask = 1'h1;
  assign mem_MPORT_228_en = reset;
  assign mem_MPORT_229_data = 32'h0;
  assign mem_MPORT_229_addr = 8'he5;
  assign mem_MPORT_229_mask = 1'h1;
  assign mem_MPORT_229_en = reset;
  assign mem_MPORT_230_data = 32'h0;
  assign mem_MPORT_230_addr = 8'he6;
  assign mem_MPORT_230_mask = 1'h1;
  assign mem_MPORT_230_en = reset;
  assign mem_MPORT_231_data = 32'h0;
  assign mem_MPORT_231_addr = 8'he7;
  assign mem_MPORT_231_mask = 1'h1;
  assign mem_MPORT_231_en = reset;
  assign mem_MPORT_232_data = 32'h0;
  assign mem_MPORT_232_addr = 8'he8;
  assign mem_MPORT_232_mask = 1'h1;
  assign mem_MPORT_232_en = reset;
  assign mem_MPORT_233_data = 32'h0;
  assign mem_MPORT_233_addr = 8'he9;
  assign mem_MPORT_233_mask = 1'h1;
  assign mem_MPORT_233_en = reset;
  assign mem_MPORT_234_data = 32'h0;
  assign mem_MPORT_234_addr = 8'hea;
  assign mem_MPORT_234_mask = 1'h1;
  assign mem_MPORT_234_en = reset;
  assign mem_MPORT_235_data = 32'h0;
  assign mem_MPORT_235_addr = 8'heb;
  assign mem_MPORT_235_mask = 1'h1;
  assign mem_MPORT_235_en = reset;
  assign mem_MPORT_236_data = 32'h0;
  assign mem_MPORT_236_addr = 8'hec;
  assign mem_MPORT_236_mask = 1'h1;
  assign mem_MPORT_236_en = reset;
  assign mem_MPORT_237_data = 32'h0;
  assign mem_MPORT_237_addr = 8'hed;
  assign mem_MPORT_237_mask = 1'h1;
  assign mem_MPORT_237_en = reset;
  assign mem_MPORT_238_data = 32'h0;
  assign mem_MPORT_238_addr = 8'hee;
  assign mem_MPORT_238_mask = 1'h1;
  assign mem_MPORT_238_en = reset;
  assign mem_MPORT_239_data = 32'h0;
  assign mem_MPORT_239_addr = 8'hef;
  assign mem_MPORT_239_mask = 1'h1;
  assign mem_MPORT_239_en = reset;
  assign mem_MPORT_240_data = 32'h0;
  assign mem_MPORT_240_addr = 8'hf0;
  assign mem_MPORT_240_mask = 1'h1;
  assign mem_MPORT_240_en = reset;
  assign mem_MPORT_241_data = 32'h0;
  assign mem_MPORT_241_addr = 8'hf1;
  assign mem_MPORT_241_mask = 1'h1;
  assign mem_MPORT_241_en = reset;
  assign mem_MPORT_242_data = 32'h0;
  assign mem_MPORT_242_addr = 8'hf2;
  assign mem_MPORT_242_mask = 1'h1;
  assign mem_MPORT_242_en = reset;
  assign mem_MPORT_243_data = 32'h0;
  assign mem_MPORT_243_addr = 8'hf3;
  assign mem_MPORT_243_mask = 1'h1;
  assign mem_MPORT_243_en = reset;
  assign mem_MPORT_244_data = 32'h0;
  assign mem_MPORT_244_addr = 8'hf4;
  assign mem_MPORT_244_mask = 1'h1;
  assign mem_MPORT_244_en = reset;
  assign mem_MPORT_245_data = 32'h0;
  assign mem_MPORT_245_addr = 8'hf5;
  assign mem_MPORT_245_mask = 1'h1;
  assign mem_MPORT_245_en = reset;
  assign mem_MPORT_246_data = 32'h0;
  assign mem_MPORT_246_addr = 8'hf6;
  assign mem_MPORT_246_mask = 1'h1;
  assign mem_MPORT_246_en = reset;
  assign mem_MPORT_247_data = 32'h0;
  assign mem_MPORT_247_addr = 8'hf7;
  assign mem_MPORT_247_mask = 1'h1;
  assign mem_MPORT_247_en = reset;
  assign mem_MPORT_248_data = 32'h0;
  assign mem_MPORT_248_addr = 8'hf8;
  assign mem_MPORT_248_mask = 1'h1;
  assign mem_MPORT_248_en = reset;
  assign mem_MPORT_249_data = 32'h0;
  assign mem_MPORT_249_addr = 8'hf9;
  assign mem_MPORT_249_mask = 1'h1;
  assign mem_MPORT_249_en = reset;
  assign mem_MPORT_250_data = 32'h0;
  assign mem_MPORT_250_addr = 8'hfa;
  assign mem_MPORT_250_mask = 1'h1;
  assign mem_MPORT_250_en = reset;
  assign mem_MPORT_251_data = 32'h0;
  assign mem_MPORT_251_addr = 8'hfb;
  assign mem_MPORT_251_mask = 1'h1;
  assign mem_MPORT_251_en = reset;
  assign mem_MPORT_252_data = 32'h0;
  assign mem_MPORT_252_addr = 8'hfc;
  assign mem_MPORT_252_mask = 1'h1;
  assign mem_MPORT_252_en = reset;
  assign mem_MPORT_253_data = 32'h0;
  assign mem_MPORT_253_addr = 8'hfd;
  assign mem_MPORT_253_mask = 1'h1;
  assign mem_MPORT_253_en = reset;
  assign mem_MPORT_254_data = 32'h0;
  assign mem_MPORT_254_addr = 8'hfe;
  assign mem_MPORT_254_mask = 1'h1;
  assign mem_MPORT_254_en = reset;
  assign mem_MPORT_255_data = 32'h0;
  assign mem_MPORT_255_addr = 8'hff;
  assign mem_MPORT_255_mask = 1'h1;
  assign mem_MPORT_255_en = reset;
  assign mem_MPORT_256_data = io_w_data;
  assign mem_MPORT_256_addr = io_w_addr;
  assign mem_MPORT_256_mask = 1'h1;
  assign mem_MPORT_256_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_129_en & mem_MPORT_129_mask) begin
      mem[mem_MPORT_129_addr] <= mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_130_en & mem_MPORT_130_mask) begin
      mem[mem_MPORT_130_addr] <= mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_131_en & mem_MPORT_131_mask) begin
      mem[mem_MPORT_131_addr] <= mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_132_en & mem_MPORT_132_mask) begin
      mem[mem_MPORT_132_addr] <= mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_133_en & mem_MPORT_133_mask) begin
      mem[mem_MPORT_133_addr] <= mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_134_en & mem_MPORT_134_mask) begin
      mem[mem_MPORT_134_addr] <= mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_135_en & mem_MPORT_135_mask) begin
      mem[mem_MPORT_135_addr] <= mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_136_en & mem_MPORT_136_mask) begin
      mem[mem_MPORT_136_addr] <= mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_137_en & mem_MPORT_137_mask) begin
      mem[mem_MPORT_137_addr] <= mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_138_en & mem_MPORT_138_mask) begin
      mem[mem_MPORT_138_addr] <= mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_139_en & mem_MPORT_139_mask) begin
      mem[mem_MPORT_139_addr] <= mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_140_en & mem_MPORT_140_mask) begin
      mem[mem_MPORT_140_addr] <= mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_141_en & mem_MPORT_141_mask) begin
      mem[mem_MPORT_141_addr] <= mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_142_en & mem_MPORT_142_mask) begin
      mem[mem_MPORT_142_addr] <= mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_143_en & mem_MPORT_143_mask) begin
      mem[mem_MPORT_143_addr] <= mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_144_en & mem_MPORT_144_mask) begin
      mem[mem_MPORT_144_addr] <= mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_145_en & mem_MPORT_145_mask) begin
      mem[mem_MPORT_145_addr] <= mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_146_en & mem_MPORT_146_mask) begin
      mem[mem_MPORT_146_addr] <= mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_147_en & mem_MPORT_147_mask) begin
      mem[mem_MPORT_147_addr] <= mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_148_en & mem_MPORT_148_mask) begin
      mem[mem_MPORT_148_addr] <= mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_149_en & mem_MPORT_149_mask) begin
      mem[mem_MPORT_149_addr] <= mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_150_en & mem_MPORT_150_mask) begin
      mem[mem_MPORT_150_addr] <= mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_151_en & mem_MPORT_151_mask) begin
      mem[mem_MPORT_151_addr] <= mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_152_en & mem_MPORT_152_mask) begin
      mem[mem_MPORT_152_addr] <= mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_153_en & mem_MPORT_153_mask) begin
      mem[mem_MPORT_153_addr] <= mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_154_en & mem_MPORT_154_mask) begin
      mem[mem_MPORT_154_addr] <= mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_155_en & mem_MPORT_155_mask) begin
      mem[mem_MPORT_155_addr] <= mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_156_en & mem_MPORT_156_mask) begin
      mem[mem_MPORT_156_addr] <= mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_157_en & mem_MPORT_157_mask) begin
      mem[mem_MPORT_157_addr] <= mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_158_en & mem_MPORT_158_mask) begin
      mem[mem_MPORT_158_addr] <= mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_159_en & mem_MPORT_159_mask) begin
      mem[mem_MPORT_159_addr] <= mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_160_en & mem_MPORT_160_mask) begin
      mem[mem_MPORT_160_addr] <= mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_161_en & mem_MPORT_161_mask) begin
      mem[mem_MPORT_161_addr] <= mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_162_en & mem_MPORT_162_mask) begin
      mem[mem_MPORT_162_addr] <= mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_163_en & mem_MPORT_163_mask) begin
      mem[mem_MPORT_163_addr] <= mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_164_en & mem_MPORT_164_mask) begin
      mem[mem_MPORT_164_addr] <= mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_165_en & mem_MPORT_165_mask) begin
      mem[mem_MPORT_165_addr] <= mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_166_en & mem_MPORT_166_mask) begin
      mem[mem_MPORT_166_addr] <= mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_167_en & mem_MPORT_167_mask) begin
      mem[mem_MPORT_167_addr] <= mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_168_en & mem_MPORT_168_mask) begin
      mem[mem_MPORT_168_addr] <= mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_169_en & mem_MPORT_169_mask) begin
      mem[mem_MPORT_169_addr] <= mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_170_en & mem_MPORT_170_mask) begin
      mem[mem_MPORT_170_addr] <= mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_171_en & mem_MPORT_171_mask) begin
      mem[mem_MPORT_171_addr] <= mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_172_en & mem_MPORT_172_mask) begin
      mem[mem_MPORT_172_addr] <= mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_173_en & mem_MPORT_173_mask) begin
      mem[mem_MPORT_173_addr] <= mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_174_en & mem_MPORT_174_mask) begin
      mem[mem_MPORT_174_addr] <= mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_175_en & mem_MPORT_175_mask) begin
      mem[mem_MPORT_175_addr] <= mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_176_en & mem_MPORT_176_mask) begin
      mem[mem_MPORT_176_addr] <= mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_177_en & mem_MPORT_177_mask) begin
      mem[mem_MPORT_177_addr] <= mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_178_en & mem_MPORT_178_mask) begin
      mem[mem_MPORT_178_addr] <= mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_179_en & mem_MPORT_179_mask) begin
      mem[mem_MPORT_179_addr] <= mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_180_en & mem_MPORT_180_mask) begin
      mem[mem_MPORT_180_addr] <= mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_181_en & mem_MPORT_181_mask) begin
      mem[mem_MPORT_181_addr] <= mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_182_en & mem_MPORT_182_mask) begin
      mem[mem_MPORT_182_addr] <= mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_183_en & mem_MPORT_183_mask) begin
      mem[mem_MPORT_183_addr] <= mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_184_en & mem_MPORT_184_mask) begin
      mem[mem_MPORT_184_addr] <= mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_185_en & mem_MPORT_185_mask) begin
      mem[mem_MPORT_185_addr] <= mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_186_en & mem_MPORT_186_mask) begin
      mem[mem_MPORT_186_addr] <= mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_187_en & mem_MPORT_187_mask) begin
      mem[mem_MPORT_187_addr] <= mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_188_en & mem_MPORT_188_mask) begin
      mem[mem_MPORT_188_addr] <= mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_189_en & mem_MPORT_189_mask) begin
      mem[mem_MPORT_189_addr] <= mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_190_en & mem_MPORT_190_mask) begin
      mem[mem_MPORT_190_addr] <= mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_191_en & mem_MPORT_191_mask) begin
      mem[mem_MPORT_191_addr] <= mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_192_en & mem_MPORT_192_mask) begin
      mem[mem_MPORT_192_addr] <= mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_193_en & mem_MPORT_193_mask) begin
      mem[mem_MPORT_193_addr] <= mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_194_en & mem_MPORT_194_mask) begin
      mem[mem_MPORT_194_addr] <= mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_195_en & mem_MPORT_195_mask) begin
      mem[mem_MPORT_195_addr] <= mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_196_en & mem_MPORT_196_mask) begin
      mem[mem_MPORT_196_addr] <= mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_197_en & mem_MPORT_197_mask) begin
      mem[mem_MPORT_197_addr] <= mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_198_en & mem_MPORT_198_mask) begin
      mem[mem_MPORT_198_addr] <= mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_199_en & mem_MPORT_199_mask) begin
      mem[mem_MPORT_199_addr] <= mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_200_en & mem_MPORT_200_mask) begin
      mem[mem_MPORT_200_addr] <= mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_201_en & mem_MPORT_201_mask) begin
      mem[mem_MPORT_201_addr] <= mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_202_en & mem_MPORT_202_mask) begin
      mem[mem_MPORT_202_addr] <= mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_203_en & mem_MPORT_203_mask) begin
      mem[mem_MPORT_203_addr] <= mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_204_en & mem_MPORT_204_mask) begin
      mem[mem_MPORT_204_addr] <= mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_205_en & mem_MPORT_205_mask) begin
      mem[mem_MPORT_205_addr] <= mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_206_en & mem_MPORT_206_mask) begin
      mem[mem_MPORT_206_addr] <= mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_207_en & mem_MPORT_207_mask) begin
      mem[mem_MPORT_207_addr] <= mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_208_en & mem_MPORT_208_mask) begin
      mem[mem_MPORT_208_addr] <= mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_209_en & mem_MPORT_209_mask) begin
      mem[mem_MPORT_209_addr] <= mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_210_en & mem_MPORT_210_mask) begin
      mem[mem_MPORT_210_addr] <= mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_211_en & mem_MPORT_211_mask) begin
      mem[mem_MPORT_211_addr] <= mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_212_en & mem_MPORT_212_mask) begin
      mem[mem_MPORT_212_addr] <= mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_213_en & mem_MPORT_213_mask) begin
      mem[mem_MPORT_213_addr] <= mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_214_en & mem_MPORT_214_mask) begin
      mem[mem_MPORT_214_addr] <= mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_215_en & mem_MPORT_215_mask) begin
      mem[mem_MPORT_215_addr] <= mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_216_en & mem_MPORT_216_mask) begin
      mem[mem_MPORT_216_addr] <= mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_217_en & mem_MPORT_217_mask) begin
      mem[mem_MPORT_217_addr] <= mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_218_en & mem_MPORT_218_mask) begin
      mem[mem_MPORT_218_addr] <= mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_219_en & mem_MPORT_219_mask) begin
      mem[mem_MPORT_219_addr] <= mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_220_en & mem_MPORT_220_mask) begin
      mem[mem_MPORT_220_addr] <= mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_221_en & mem_MPORT_221_mask) begin
      mem[mem_MPORT_221_addr] <= mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_222_en & mem_MPORT_222_mask) begin
      mem[mem_MPORT_222_addr] <= mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_223_en & mem_MPORT_223_mask) begin
      mem[mem_MPORT_223_addr] <= mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_224_en & mem_MPORT_224_mask) begin
      mem[mem_MPORT_224_addr] <= mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_225_en & mem_MPORT_225_mask) begin
      mem[mem_MPORT_225_addr] <= mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_226_en & mem_MPORT_226_mask) begin
      mem[mem_MPORT_226_addr] <= mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_227_en & mem_MPORT_227_mask) begin
      mem[mem_MPORT_227_addr] <= mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_228_en & mem_MPORT_228_mask) begin
      mem[mem_MPORT_228_addr] <= mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_229_en & mem_MPORT_229_mask) begin
      mem[mem_MPORT_229_addr] <= mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_230_en & mem_MPORT_230_mask) begin
      mem[mem_MPORT_230_addr] <= mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_231_en & mem_MPORT_231_mask) begin
      mem[mem_MPORT_231_addr] <= mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_232_en & mem_MPORT_232_mask) begin
      mem[mem_MPORT_232_addr] <= mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_233_en & mem_MPORT_233_mask) begin
      mem[mem_MPORT_233_addr] <= mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_234_en & mem_MPORT_234_mask) begin
      mem[mem_MPORT_234_addr] <= mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_235_en & mem_MPORT_235_mask) begin
      mem[mem_MPORT_235_addr] <= mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_236_en & mem_MPORT_236_mask) begin
      mem[mem_MPORT_236_addr] <= mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_237_en & mem_MPORT_237_mask) begin
      mem[mem_MPORT_237_addr] <= mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_238_en & mem_MPORT_238_mask) begin
      mem[mem_MPORT_238_addr] <= mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_239_en & mem_MPORT_239_mask) begin
      mem[mem_MPORT_239_addr] <= mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_240_en & mem_MPORT_240_mask) begin
      mem[mem_MPORT_240_addr] <= mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_241_en & mem_MPORT_241_mask) begin
      mem[mem_MPORT_241_addr] <= mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_242_en & mem_MPORT_242_mask) begin
      mem[mem_MPORT_242_addr] <= mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_243_en & mem_MPORT_243_mask) begin
      mem[mem_MPORT_243_addr] <= mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_244_en & mem_MPORT_244_mask) begin
      mem[mem_MPORT_244_addr] <= mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_245_en & mem_MPORT_245_mask) begin
      mem[mem_MPORT_245_addr] <= mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_246_en & mem_MPORT_246_mask) begin
      mem[mem_MPORT_246_addr] <= mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_247_en & mem_MPORT_247_mask) begin
      mem[mem_MPORT_247_addr] <= mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_248_en & mem_MPORT_248_mask) begin
      mem[mem_MPORT_248_addr] <= mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_249_en & mem_MPORT_249_mask) begin
      mem[mem_MPORT_249_addr] <= mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_250_en & mem_MPORT_250_mask) begin
      mem[mem_MPORT_250_addr] <= mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_251_en & mem_MPORT_251_mask) begin
      mem[mem_MPORT_251_addr] <= mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_252_en & mem_MPORT_252_mask) begin
      mem[mem_MPORT_252_addr] <= mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_253_en & mem_MPORT_253_mask) begin
      mem[mem_MPORT_253_addr] <= mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_254_en & mem_MPORT_254_mask) begin
      mem[mem_MPORT_254_addr] <= mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_255_en & mem_MPORT_255_mask) begin
      mem[mem_MPORT_255_addr] <= mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_256_en & mem_MPORT_256_mask) begin
      mem[mem_MPORT_256_addr] <= mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_10(
  input         clock,
  input         reset,
  input  [7:0]  io_r_addr,
  output [31:0] io_r_data_0,
  output [31:0] io_r_data_1,
  output [31:0] io_r_data_2,
  output [31:0] io_r_data_3,
  input         io_w_en,
  input  [7:0]  io_w_addr,
  input  [31:0] io_w_data_0,
  input  [31:0] io_w_data_1,
  input  [31:0] io_w_data_2,
  input  [31:0] io_w_data_3,
  input  [3:0]  io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [31:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P_80 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P_80 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P_80 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P_80 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
endmodule
module DataBankArray_1(
  input         clock,
  input         reset,
  output        io_read_req_ready,
  input         io_read_req_valid,
  input  [7:0]  io_read_req_bits_set,
  output [31:0] io_read_resp_0_0,
  output [31:0] io_read_resp_0_1,
  output [31:0] io_read_resp_0_2,
  output [31:0] io_read_resp_0_3,
  output [31:0] io_read_resp_1_0,
  output [31:0] io_read_resp_1_1,
  output [31:0] io_read_resp_1_2,
  output [31:0] io_read_resp_1_3,
  output [31:0] io_read_resp_2_0,
  output [31:0] io_read_resp_2_1,
  output [31:0] io_read_resp_2_2,
  output [31:0] io_read_resp_2_3,
  output [31:0] io_read_resp_3_0,
  output [31:0] io_read_resp_3_1,
  output [31:0] io_read_resp_3_2,
  output [31:0] io_read_resp_3_3,
  output [31:0] io_read_resp_4_0,
  output [31:0] io_read_resp_4_1,
  output [31:0] io_read_resp_4_2,
  output [31:0] io_read_resp_4_3,
  output [31:0] io_read_resp_5_0,
  output [31:0] io_read_resp_5_1,
  output [31:0] io_read_resp_5_2,
  output [31:0] io_read_resp_5_3,
  output [31:0] io_read_resp_6_0,
  output [31:0] io_read_resp_6_1,
  output [31:0] io_read_resp_6_2,
  output [31:0] io_read_resp_6_3,
  output [31:0] io_read_resp_7_0,
  output [31:0] io_read_resp_7_1,
  output [31:0] io_read_resp_7_2,
  output [31:0] io_read_resp_7_3,
  output        io_write_req_ready,
  input         io_write_req_valid,
  input  [7:0]  io_write_req_bits_set,
  input  [31:0] io_write_req_bits_data_0,
  input  [31:0] io_write_req_bits_data_1,
  input  [31:0] io_write_req_bits_data_2,
  input  [31:0] io_write_req_bits_data_3,
  input  [3:0]  io_write_req_bits_blockMask,
  input  [7:0]  io_write_req_bits_way
);
  wire  dataBanks_0_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_0_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_0_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_0_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_0_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_0_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_0_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_1_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_1_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_1_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_1_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_1_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_2_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_2_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_2_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_2_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_2_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_3_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_3_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_3_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_3_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_3_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_4_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_4_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_4_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_4_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_4_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_4_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_4_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_5_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_5_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_5_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_5_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_5_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_5_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_5_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_6_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_6_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_6_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_6_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_6_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_6_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_6_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  dataBanks_7_clock; // @[SRAM_1.scala 255:31]
  wire  dataBanks_7_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_7_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire  dataBanks_7_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] dataBanks_7_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [31:0] dataBanks_7_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [3:0] dataBanks_7_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  ren = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  wire  _wen_T_1 = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  SRAMArray_2P_10 dataBanks_0 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_0_clock),
    .reset(dataBanks_0_reset),
    .io_r_addr(dataBanks_0_io_r_addr),
    .io_r_data_0(dataBanks_0_io_r_data_0),
    .io_r_data_1(dataBanks_0_io_r_data_1),
    .io_r_data_2(dataBanks_0_io_r_data_2),
    .io_r_data_3(dataBanks_0_io_r_data_3),
    .io_w_en(dataBanks_0_io_w_en),
    .io_w_addr(dataBanks_0_io_w_addr),
    .io_w_data_0(dataBanks_0_io_w_data_0),
    .io_w_data_1(dataBanks_0_io_w_data_1),
    .io_w_data_2(dataBanks_0_io_w_data_2),
    .io_w_data_3(dataBanks_0_io_w_data_3),
    .io_w_maskOH(dataBanks_0_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_1 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_1_clock),
    .reset(dataBanks_1_reset),
    .io_r_addr(dataBanks_1_io_r_addr),
    .io_r_data_0(dataBanks_1_io_r_data_0),
    .io_r_data_1(dataBanks_1_io_r_data_1),
    .io_r_data_2(dataBanks_1_io_r_data_2),
    .io_r_data_3(dataBanks_1_io_r_data_3),
    .io_w_en(dataBanks_1_io_w_en),
    .io_w_addr(dataBanks_1_io_w_addr),
    .io_w_data_0(dataBanks_1_io_w_data_0),
    .io_w_data_1(dataBanks_1_io_w_data_1),
    .io_w_data_2(dataBanks_1_io_w_data_2),
    .io_w_data_3(dataBanks_1_io_w_data_3),
    .io_w_maskOH(dataBanks_1_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_2 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_2_clock),
    .reset(dataBanks_2_reset),
    .io_r_addr(dataBanks_2_io_r_addr),
    .io_r_data_0(dataBanks_2_io_r_data_0),
    .io_r_data_1(dataBanks_2_io_r_data_1),
    .io_r_data_2(dataBanks_2_io_r_data_2),
    .io_r_data_3(dataBanks_2_io_r_data_3),
    .io_w_en(dataBanks_2_io_w_en),
    .io_w_addr(dataBanks_2_io_w_addr),
    .io_w_data_0(dataBanks_2_io_w_data_0),
    .io_w_data_1(dataBanks_2_io_w_data_1),
    .io_w_data_2(dataBanks_2_io_w_data_2),
    .io_w_data_3(dataBanks_2_io_w_data_3),
    .io_w_maskOH(dataBanks_2_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_3 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_3_clock),
    .reset(dataBanks_3_reset),
    .io_r_addr(dataBanks_3_io_r_addr),
    .io_r_data_0(dataBanks_3_io_r_data_0),
    .io_r_data_1(dataBanks_3_io_r_data_1),
    .io_r_data_2(dataBanks_3_io_r_data_2),
    .io_r_data_3(dataBanks_3_io_r_data_3),
    .io_w_en(dataBanks_3_io_w_en),
    .io_w_addr(dataBanks_3_io_w_addr),
    .io_w_data_0(dataBanks_3_io_w_data_0),
    .io_w_data_1(dataBanks_3_io_w_data_1),
    .io_w_data_2(dataBanks_3_io_w_data_2),
    .io_w_data_3(dataBanks_3_io_w_data_3),
    .io_w_maskOH(dataBanks_3_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_4 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_4_clock),
    .reset(dataBanks_4_reset),
    .io_r_addr(dataBanks_4_io_r_addr),
    .io_r_data_0(dataBanks_4_io_r_data_0),
    .io_r_data_1(dataBanks_4_io_r_data_1),
    .io_r_data_2(dataBanks_4_io_r_data_2),
    .io_r_data_3(dataBanks_4_io_r_data_3),
    .io_w_en(dataBanks_4_io_w_en),
    .io_w_addr(dataBanks_4_io_w_addr),
    .io_w_data_0(dataBanks_4_io_w_data_0),
    .io_w_data_1(dataBanks_4_io_w_data_1),
    .io_w_data_2(dataBanks_4_io_w_data_2),
    .io_w_data_3(dataBanks_4_io_w_data_3),
    .io_w_maskOH(dataBanks_4_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_5 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_5_clock),
    .reset(dataBanks_5_reset),
    .io_r_addr(dataBanks_5_io_r_addr),
    .io_r_data_0(dataBanks_5_io_r_data_0),
    .io_r_data_1(dataBanks_5_io_r_data_1),
    .io_r_data_2(dataBanks_5_io_r_data_2),
    .io_r_data_3(dataBanks_5_io_r_data_3),
    .io_w_en(dataBanks_5_io_w_en),
    .io_w_addr(dataBanks_5_io_w_addr),
    .io_w_data_0(dataBanks_5_io_w_data_0),
    .io_w_data_1(dataBanks_5_io_w_data_1),
    .io_w_data_2(dataBanks_5_io_w_data_2),
    .io_w_data_3(dataBanks_5_io_w_data_3),
    .io_w_maskOH(dataBanks_5_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_6 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_6_clock),
    .reset(dataBanks_6_reset),
    .io_r_addr(dataBanks_6_io_r_addr),
    .io_r_data_0(dataBanks_6_io_r_data_0),
    .io_r_data_1(dataBanks_6_io_r_data_1),
    .io_r_data_2(dataBanks_6_io_r_data_2),
    .io_r_data_3(dataBanks_6_io_r_data_3),
    .io_w_en(dataBanks_6_io_w_en),
    .io_w_addr(dataBanks_6_io_w_addr),
    .io_w_data_0(dataBanks_6_io_w_data_0),
    .io_w_data_1(dataBanks_6_io_w_data_1),
    .io_w_data_2(dataBanks_6_io_w_data_2),
    .io_w_data_3(dataBanks_6_io_w_data_3),
    .io_w_maskOH(dataBanks_6_io_w_maskOH)
  );
  SRAMArray_2P_10 dataBanks_7 ( // @[SRAM_1.scala 255:31]
    .clock(dataBanks_7_clock),
    .reset(dataBanks_7_reset),
    .io_r_addr(dataBanks_7_io_r_addr),
    .io_r_data_0(dataBanks_7_io_r_data_0),
    .io_r_data_1(dataBanks_7_io_r_data_1),
    .io_r_data_2(dataBanks_7_io_r_data_2),
    .io_r_data_3(dataBanks_7_io_r_data_3),
    .io_w_en(dataBanks_7_io_w_en),
    .io_w_addr(dataBanks_7_io_w_addr),
    .io_w_data_0(dataBanks_7_io_w_data_0),
    .io_w_data_1(dataBanks_7_io_w_data_1),
    .io_w_data_2(dataBanks_7_io_w_data_2),
    .io_w_data_3(dataBanks_7_io_w_data_3),
    .io_w_maskOH(dataBanks_7_io_w_maskOH)
  );
  assign io_read_req_ready = 1'h1; // @[DataBank.scala 46:23]
  assign io_read_resp_0_0 = ren ? dataBanks_0_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_1 = ren ? dataBanks_0_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_2 = ren ? dataBanks_0_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_0_3 = ren ? dataBanks_0_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_0 = ren ? dataBanks_1_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_1 = ren ? dataBanks_1_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_2 = ren ? dataBanks_1_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_1_3 = ren ? dataBanks_1_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_0 = ren ? dataBanks_2_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_1 = ren ? dataBanks_2_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_2 = ren ? dataBanks_2_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_2_3 = ren ? dataBanks_2_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_0 = ren ? dataBanks_3_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_1 = ren ? dataBanks_3_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_2 = ren ? dataBanks_3_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_3_3 = ren ? dataBanks_3_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_0 = ren ? dataBanks_4_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_1 = ren ? dataBanks_4_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_2 = ren ? dataBanks_4_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_4_3 = ren ? dataBanks_4_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_0 = ren ? dataBanks_5_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_1 = ren ? dataBanks_5_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_2 = ren ? dataBanks_5_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_5_3 = ren ? dataBanks_5_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_0 = ren ? dataBanks_6_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_1 = ren ? dataBanks_6_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_2 = ren ? dataBanks_6_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_6_3 = ren ? dataBanks_6_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_0 = ren ? dataBanks_7_io_r_data_0 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_1 = ren ? dataBanks_7_io_r_data_1 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_2 = ren ? dataBanks_7_io_r_data_2 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_7_3 = ren ? dataBanks_7_io_r_data_3 : 32'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_write_req_ready = 1'h1; // @[DataBank.scala 55:28]
  assign dataBanks_0_clock = clock;
  assign dataBanks_0_reset = reset;
  assign dataBanks_0_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_0_io_w_en = io_write_req_bits_way[0] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_0_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_0_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_0_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_1_clock = clock;
  assign dataBanks_1_reset = reset;
  assign dataBanks_1_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_1_io_w_en = io_write_req_bits_way[1] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_1_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_1_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_1_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_2_clock = clock;
  assign dataBanks_2_reset = reset;
  assign dataBanks_2_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_2_io_w_en = io_write_req_bits_way[2] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_2_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_2_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_2_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_3_clock = clock;
  assign dataBanks_3_reset = reset;
  assign dataBanks_3_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_3_io_w_en = io_write_req_bits_way[3] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_3_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_3_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_3_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_4_clock = clock;
  assign dataBanks_4_reset = reset;
  assign dataBanks_4_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_4_io_w_en = io_write_req_bits_way[4] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_4_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_4_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_4_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_5_clock = clock;
  assign dataBanks_5_reset = reset;
  assign dataBanks_5_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_5_io_w_en = io_write_req_bits_way[5] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_5_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_5_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_5_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_6_clock = clock;
  assign dataBanks_6_reset = reset;
  assign dataBanks_6_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_6_io_w_en = io_write_req_bits_way[6] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_6_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_6_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_6_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
  assign dataBanks_7_clock = clock;
  assign dataBanks_7_reset = reset;
  assign dataBanks_7_io_r_addr = io_read_req_bits_set; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign dataBanks_7_io_w_en = io_write_req_bits_way[7] & _wen_T_1; // @[DataBank.scala 53:44]
  assign dataBanks_7_io_w_addr = io_write_req_bits_set; // @[DataBank.scala 56:19 SRAM_1.scala 222:19]
  assign dataBanks_7_io_w_data_0 = io_write_req_bits_data_0; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_1 = io_write_req_bits_data_1; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_2 = io_write_req_bits_data_2; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_data_3 = io_write_req_bits_data_3; // @[DataBank.scala 56:19 SRAM_1.scala 223:19]
  assign dataBanks_7_io_w_maskOH = io_write_req_bits_blockMask; // @[DataBank.scala 56:19 SRAM_1.scala 224:21]
endmodule
module BankRAM_2P_112(
  input         clock,
  input         reset,
  input  [7:0]  io_r_addr,
  output [19:0] io_r_data,
  input         io_w_en,
  input  [7:0]  io_w_addr,
  input  [19:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] mem [0:255]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_129_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_130_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_131_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_132_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_133_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_134_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_135_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_136_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_137_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_138_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_139_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_140_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_141_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_142_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_143_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_144_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_145_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_146_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_147_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_148_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_149_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_150_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_151_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_152_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_153_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_154_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_155_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_156_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_157_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_158_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_159_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_160_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_161_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_162_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_163_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_164_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_165_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_166_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_167_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_168_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_169_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_170_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_171_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_172_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_173_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_174_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_175_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_176_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_177_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_178_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_179_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_180_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_181_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_182_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_183_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_184_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_185_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_186_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_187_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_188_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_189_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_190_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_191_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_192_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_193_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_194_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_195_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_196_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_197_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_198_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_199_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_200_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_201_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_202_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_203_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_204_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_205_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_206_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_207_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_208_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_209_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_210_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_211_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_212_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_213_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_214_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_215_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_216_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_217_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_218_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_219_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_220_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_221_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_222_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_223_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_224_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_225_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_226_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_227_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_228_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_229_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_230_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_231_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_232_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_233_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_234_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_235_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_236_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_237_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_238_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_239_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_240_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_241_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_242_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_243_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_244_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_245_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_246_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_247_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_248_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_249_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_250_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_251_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_252_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_253_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_254_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_255_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_en; // @[SRAM_1.scala 63:26]
  wire [19:0] mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_256_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [7:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 20'h0;
  assign mem_MPORT_addr = 8'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 20'h0;
  assign mem_MPORT_1_addr = 8'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 20'h0;
  assign mem_MPORT_2_addr = 8'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 20'h0;
  assign mem_MPORT_3_addr = 8'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 20'h0;
  assign mem_MPORT_4_addr = 8'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 20'h0;
  assign mem_MPORT_5_addr = 8'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 20'h0;
  assign mem_MPORT_6_addr = 8'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 20'h0;
  assign mem_MPORT_7_addr = 8'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 20'h0;
  assign mem_MPORT_8_addr = 8'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 20'h0;
  assign mem_MPORT_9_addr = 8'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 20'h0;
  assign mem_MPORT_10_addr = 8'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 20'h0;
  assign mem_MPORT_11_addr = 8'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 20'h0;
  assign mem_MPORT_12_addr = 8'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 20'h0;
  assign mem_MPORT_13_addr = 8'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 20'h0;
  assign mem_MPORT_14_addr = 8'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 20'h0;
  assign mem_MPORT_15_addr = 8'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 20'h0;
  assign mem_MPORT_16_addr = 8'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 20'h0;
  assign mem_MPORT_17_addr = 8'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 20'h0;
  assign mem_MPORT_18_addr = 8'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 20'h0;
  assign mem_MPORT_19_addr = 8'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 20'h0;
  assign mem_MPORT_20_addr = 8'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 20'h0;
  assign mem_MPORT_21_addr = 8'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 20'h0;
  assign mem_MPORT_22_addr = 8'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 20'h0;
  assign mem_MPORT_23_addr = 8'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 20'h0;
  assign mem_MPORT_24_addr = 8'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 20'h0;
  assign mem_MPORT_25_addr = 8'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 20'h0;
  assign mem_MPORT_26_addr = 8'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 20'h0;
  assign mem_MPORT_27_addr = 8'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 20'h0;
  assign mem_MPORT_28_addr = 8'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 20'h0;
  assign mem_MPORT_29_addr = 8'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 20'h0;
  assign mem_MPORT_30_addr = 8'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 20'h0;
  assign mem_MPORT_31_addr = 8'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 20'h0;
  assign mem_MPORT_32_addr = 8'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 20'h0;
  assign mem_MPORT_33_addr = 8'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 20'h0;
  assign mem_MPORT_34_addr = 8'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 20'h0;
  assign mem_MPORT_35_addr = 8'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 20'h0;
  assign mem_MPORT_36_addr = 8'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 20'h0;
  assign mem_MPORT_37_addr = 8'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 20'h0;
  assign mem_MPORT_38_addr = 8'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 20'h0;
  assign mem_MPORT_39_addr = 8'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 20'h0;
  assign mem_MPORT_40_addr = 8'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 20'h0;
  assign mem_MPORT_41_addr = 8'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 20'h0;
  assign mem_MPORT_42_addr = 8'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 20'h0;
  assign mem_MPORT_43_addr = 8'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 20'h0;
  assign mem_MPORT_44_addr = 8'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 20'h0;
  assign mem_MPORT_45_addr = 8'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 20'h0;
  assign mem_MPORT_46_addr = 8'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 20'h0;
  assign mem_MPORT_47_addr = 8'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 20'h0;
  assign mem_MPORT_48_addr = 8'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 20'h0;
  assign mem_MPORT_49_addr = 8'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 20'h0;
  assign mem_MPORT_50_addr = 8'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 20'h0;
  assign mem_MPORT_51_addr = 8'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 20'h0;
  assign mem_MPORT_52_addr = 8'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 20'h0;
  assign mem_MPORT_53_addr = 8'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 20'h0;
  assign mem_MPORT_54_addr = 8'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 20'h0;
  assign mem_MPORT_55_addr = 8'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 20'h0;
  assign mem_MPORT_56_addr = 8'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 20'h0;
  assign mem_MPORT_57_addr = 8'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 20'h0;
  assign mem_MPORT_58_addr = 8'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 20'h0;
  assign mem_MPORT_59_addr = 8'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 20'h0;
  assign mem_MPORT_60_addr = 8'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 20'h0;
  assign mem_MPORT_61_addr = 8'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 20'h0;
  assign mem_MPORT_62_addr = 8'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 20'h0;
  assign mem_MPORT_63_addr = 8'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 20'h0;
  assign mem_MPORT_64_addr = 8'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 20'h0;
  assign mem_MPORT_65_addr = 8'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 20'h0;
  assign mem_MPORT_66_addr = 8'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 20'h0;
  assign mem_MPORT_67_addr = 8'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 20'h0;
  assign mem_MPORT_68_addr = 8'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 20'h0;
  assign mem_MPORT_69_addr = 8'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 20'h0;
  assign mem_MPORT_70_addr = 8'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 20'h0;
  assign mem_MPORT_71_addr = 8'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 20'h0;
  assign mem_MPORT_72_addr = 8'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 20'h0;
  assign mem_MPORT_73_addr = 8'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 20'h0;
  assign mem_MPORT_74_addr = 8'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 20'h0;
  assign mem_MPORT_75_addr = 8'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 20'h0;
  assign mem_MPORT_76_addr = 8'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 20'h0;
  assign mem_MPORT_77_addr = 8'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 20'h0;
  assign mem_MPORT_78_addr = 8'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 20'h0;
  assign mem_MPORT_79_addr = 8'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 20'h0;
  assign mem_MPORT_80_addr = 8'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 20'h0;
  assign mem_MPORT_81_addr = 8'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 20'h0;
  assign mem_MPORT_82_addr = 8'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 20'h0;
  assign mem_MPORT_83_addr = 8'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 20'h0;
  assign mem_MPORT_84_addr = 8'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 20'h0;
  assign mem_MPORT_85_addr = 8'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 20'h0;
  assign mem_MPORT_86_addr = 8'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 20'h0;
  assign mem_MPORT_87_addr = 8'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 20'h0;
  assign mem_MPORT_88_addr = 8'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 20'h0;
  assign mem_MPORT_89_addr = 8'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 20'h0;
  assign mem_MPORT_90_addr = 8'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 20'h0;
  assign mem_MPORT_91_addr = 8'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 20'h0;
  assign mem_MPORT_92_addr = 8'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 20'h0;
  assign mem_MPORT_93_addr = 8'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 20'h0;
  assign mem_MPORT_94_addr = 8'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 20'h0;
  assign mem_MPORT_95_addr = 8'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 20'h0;
  assign mem_MPORT_96_addr = 8'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 20'h0;
  assign mem_MPORT_97_addr = 8'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 20'h0;
  assign mem_MPORT_98_addr = 8'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 20'h0;
  assign mem_MPORT_99_addr = 8'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 20'h0;
  assign mem_MPORT_100_addr = 8'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 20'h0;
  assign mem_MPORT_101_addr = 8'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 20'h0;
  assign mem_MPORT_102_addr = 8'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 20'h0;
  assign mem_MPORT_103_addr = 8'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 20'h0;
  assign mem_MPORT_104_addr = 8'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 20'h0;
  assign mem_MPORT_105_addr = 8'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 20'h0;
  assign mem_MPORT_106_addr = 8'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 20'h0;
  assign mem_MPORT_107_addr = 8'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 20'h0;
  assign mem_MPORT_108_addr = 8'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 20'h0;
  assign mem_MPORT_109_addr = 8'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 20'h0;
  assign mem_MPORT_110_addr = 8'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 20'h0;
  assign mem_MPORT_111_addr = 8'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 20'h0;
  assign mem_MPORT_112_addr = 8'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 20'h0;
  assign mem_MPORT_113_addr = 8'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 20'h0;
  assign mem_MPORT_114_addr = 8'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 20'h0;
  assign mem_MPORT_115_addr = 8'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 20'h0;
  assign mem_MPORT_116_addr = 8'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 20'h0;
  assign mem_MPORT_117_addr = 8'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 20'h0;
  assign mem_MPORT_118_addr = 8'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 20'h0;
  assign mem_MPORT_119_addr = 8'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 20'h0;
  assign mem_MPORT_120_addr = 8'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 20'h0;
  assign mem_MPORT_121_addr = 8'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 20'h0;
  assign mem_MPORT_122_addr = 8'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 20'h0;
  assign mem_MPORT_123_addr = 8'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 20'h0;
  assign mem_MPORT_124_addr = 8'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 20'h0;
  assign mem_MPORT_125_addr = 8'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 20'h0;
  assign mem_MPORT_126_addr = 8'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 20'h0;
  assign mem_MPORT_127_addr = 8'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 20'h0;
  assign mem_MPORT_128_addr = 8'h80;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = reset;
  assign mem_MPORT_129_data = 20'h0;
  assign mem_MPORT_129_addr = 8'h81;
  assign mem_MPORT_129_mask = 1'h1;
  assign mem_MPORT_129_en = reset;
  assign mem_MPORT_130_data = 20'h0;
  assign mem_MPORT_130_addr = 8'h82;
  assign mem_MPORT_130_mask = 1'h1;
  assign mem_MPORT_130_en = reset;
  assign mem_MPORT_131_data = 20'h0;
  assign mem_MPORT_131_addr = 8'h83;
  assign mem_MPORT_131_mask = 1'h1;
  assign mem_MPORT_131_en = reset;
  assign mem_MPORT_132_data = 20'h0;
  assign mem_MPORT_132_addr = 8'h84;
  assign mem_MPORT_132_mask = 1'h1;
  assign mem_MPORT_132_en = reset;
  assign mem_MPORT_133_data = 20'h0;
  assign mem_MPORT_133_addr = 8'h85;
  assign mem_MPORT_133_mask = 1'h1;
  assign mem_MPORT_133_en = reset;
  assign mem_MPORT_134_data = 20'h0;
  assign mem_MPORT_134_addr = 8'h86;
  assign mem_MPORT_134_mask = 1'h1;
  assign mem_MPORT_134_en = reset;
  assign mem_MPORT_135_data = 20'h0;
  assign mem_MPORT_135_addr = 8'h87;
  assign mem_MPORT_135_mask = 1'h1;
  assign mem_MPORT_135_en = reset;
  assign mem_MPORT_136_data = 20'h0;
  assign mem_MPORT_136_addr = 8'h88;
  assign mem_MPORT_136_mask = 1'h1;
  assign mem_MPORT_136_en = reset;
  assign mem_MPORT_137_data = 20'h0;
  assign mem_MPORT_137_addr = 8'h89;
  assign mem_MPORT_137_mask = 1'h1;
  assign mem_MPORT_137_en = reset;
  assign mem_MPORT_138_data = 20'h0;
  assign mem_MPORT_138_addr = 8'h8a;
  assign mem_MPORT_138_mask = 1'h1;
  assign mem_MPORT_138_en = reset;
  assign mem_MPORT_139_data = 20'h0;
  assign mem_MPORT_139_addr = 8'h8b;
  assign mem_MPORT_139_mask = 1'h1;
  assign mem_MPORT_139_en = reset;
  assign mem_MPORT_140_data = 20'h0;
  assign mem_MPORT_140_addr = 8'h8c;
  assign mem_MPORT_140_mask = 1'h1;
  assign mem_MPORT_140_en = reset;
  assign mem_MPORT_141_data = 20'h0;
  assign mem_MPORT_141_addr = 8'h8d;
  assign mem_MPORT_141_mask = 1'h1;
  assign mem_MPORT_141_en = reset;
  assign mem_MPORT_142_data = 20'h0;
  assign mem_MPORT_142_addr = 8'h8e;
  assign mem_MPORT_142_mask = 1'h1;
  assign mem_MPORT_142_en = reset;
  assign mem_MPORT_143_data = 20'h0;
  assign mem_MPORT_143_addr = 8'h8f;
  assign mem_MPORT_143_mask = 1'h1;
  assign mem_MPORT_143_en = reset;
  assign mem_MPORT_144_data = 20'h0;
  assign mem_MPORT_144_addr = 8'h90;
  assign mem_MPORT_144_mask = 1'h1;
  assign mem_MPORT_144_en = reset;
  assign mem_MPORT_145_data = 20'h0;
  assign mem_MPORT_145_addr = 8'h91;
  assign mem_MPORT_145_mask = 1'h1;
  assign mem_MPORT_145_en = reset;
  assign mem_MPORT_146_data = 20'h0;
  assign mem_MPORT_146_addr = 8'h92;
  assign mem_MPORT_146_mask = 1'h1;
  assign mem_MPORT_146_en = reset;
  assign mem_MPORT_147_data = 20'h0;
  assign mem_MPORT_147_addr = 8'h93;
  assign mem_MPORT_147_mask = 1'h1;
  assign mem_MPORT_147_en = reset;
  assign mem_MPORT_148_data = 20'h0;
  assign mem_MPORT_148_addr = 8'h94;
  assign mem_MPORT_148_mask = 1'h1;
  assign mem_MPORT_148_en = reset;
  assign mem_MPORT_149_data = 20'h0;
  assign mem_MPORT_149_addr = 8'h95;
  assign mem_MPORT_149_mask = 1'h1;
  assign mem_MPORT_149_en = reset;
  assign mem_MPORT_150_data = 20'h0;
  assign mem_MPORT_150_addr = 8'h96;
  assign mem_MPORT_150_mask = 1'h1;
  assign mem_MPORT_150_en = reset;
  assign mem_MPORT_151_data = 20'h0;
  assign mem_MPORT_151_addr = 8'h97;
  assign mem_MPORT_151_mask = 1'h1;
  assign mem_MPORT_151_en = reset;
  assign mem_MPORT_152_data = 20'h0;
  assign mem_MPORT_152_addr = 8'h98;
  assign mem_MPORT_152_mask = 1'h1;
  assign mem_MPORT_152_en = reset;
  assign mem_MPORT_153_data = 20'h0;
  assign mem_MPORT_153_addr = 8'h99;
  assign mem_MPORT_153_mask = 1'h1;
  assign mem_MPORT_153_en = reset;
  assign mem_MPORT_154_data = 20'h0;
  assign mem_MPORT_154_addr = 8'h9a;
  assign mem_MPORT_154_mask = 1'h1;
  assign mem_MPORT_154_en = reset;
  assign mem_MPORT_155_data = 20'h0;
  assign mem_MPORT_155_addr = 8'h9b;
  assign mem_MPORT_155_mask = 1'h1;
  assign mem_MPORT_155_en = reset;
  assign mem_MPORT_156_data = 20'h0;
  assign mem_MPORT_156_addr = 8'h9c;
  assign mem_MPORT_156_mask = 1'h1;
  assign mem_MPORT_156_en = reset;
  assign mem_MPORT_157_data = 20'h0;
  assign mem_MPORT_157_addr = 8'h9d;
  assign mem_MPORT_157_mask = 1'h1;
  assign mem_MPORT_157_en = reset;
  assign mem_MPORT_158_data = 20'h0;
  assign mem_MPORT_158_addr = 8'h9e;
  assign mem_MPORT_158_mask = 1'h1;
  assign mem_MPORT_158_en = reset;
  assign mem_MPORT_159_data = 20'h0;
  assign mem_MPORT_159_addr = 8'h9f;
  assign mem_MPORT_159_mask = 1'h1;
  assign mem_MPORT_159_en = reset;
  assign mem_MPORT_160_data = 20'h0;
  assign mem_MPORT_160_addr = 8'ha0;
  assign mem_MPORT_160_mask = 1'h1;
  assign mem_MPORT_160_en = reset;
  assign mem_MPORT_161_data = 20'h0;
  assign mem_MPORT_161_addr = 8'ha1;
  assign mem_MPORT_161_mask = 1'h1;
  assign mem_MPORT_161_en = reset;
  assign mem_MPORT_162_data = 20'h0;
  assign mem_MPORT_162_addr = 8'ha2;
  assign mem_MPORT_162_mask = 1'h1;
  assign mem_MPORT_162_en = reset;
  assign mem_MPORT_163_data = 20'h0;
  assign mem_MPORT_163_addr = 8'ha3;
  assign mem_MPORT_163_mask = 1'h1;
  assign mem_MPORT_163_en = reset;
  assign mem_MPORT_164_data = 20'h0;
  assign mem_MPORT_164_addr = 8'ha4;
  assign mem_MPORT_164_mask = 1'h1;
  assign mem_MPORT_164_en = reset;
  assign mem_MPORT_165_data = 20'h0;
  assign mem_MPORT_165_addr = 8'ha5;
  assign mem_MPORT_165_mask = 1'h1;
  assign mem_MPORT_165_en = reset;
  assign mem_MPORT_166_data = 20'h0;
  assign mem_MPORT_166_addr = 8'ha6;
  assign mem_MPORT_166_mask = 1'h1;
  assign mem_MPORT_166_en = reset;
  assign mem_MPORT_167_data = 20'h0;
  assign mem_MPORT_167_addr = 8'ha7;
  assign mem_MPORT_167_mask = 1'h1;
  assign mem_MPORT_167_en = reset;
  assign mem_MPORT_168_data = 20'h0;
  assign mem_MPORT_168_addr = 8'ha8;
  assign mem_MPORT_168_mask = 1'h1;
  assign mem_MPORT_168_en = reset;
  assign mem_MPORT_169_data = 20'h0;
  assign mem_MPORT_169_addr = 8'ha9;
  assign mem_MPORT_169_mask = 1'h1;
  assign mem_MPORT_169_en = reset;
  assign mem_MPORT_170_data = 20'h0;
  assign mem_MPORT_170_addr = 8'haa;
  assign mem_MPORT_170_mask = 1'h1;
  assign mem_MPORT_170_en = reset;
  assign mem_MPORT_171_data = 20'h0;
  assign mem_MPORT_171_addr = 8'hab;
  assign mem_MPORT_171_mask = 1'h1;
  assign mem_MPORT_171_en = reset;
  assign mem_MPORT_172_data = 20'h0;
  assign mem_MPORT_172_addr = 8'hac;
  assign mem_MPORT_172_mask = 1'h1;
  assign mem_MPORT_172_en = reset;
  assign mem_MPORT_173_data = 20'h0;
  assign mem_MPORT_173_addr = 8'had;
  assign mem_MPORT_173_mask = 1'h1;
  assign mem_MPORT_173_en = reset;
  assign mem_MPORT_174_data = 20'h0;
  assign mem_MPORT_174_addr = 8'hae;
  assign mem_MPORT_174_mask = 1'h1;
  assign mem_MPORT_174_en = reset;
  assign mem_MPORT_175_data = 20'h0;
  assign mem_MPORT_175_addr = 8'haf;
  assign mem_MPORT_175_mask = 1'h1;
  assign mem_MPORT_175_en = reset;
  assign mem_MPORT_176_data = 20'h0;
  assign mem_MPORT_176_addr = 8'hb0;
  assign mem_MPORT_176_mask = 1'h1;
  assign mem_MPORT_176_en = reset;
  assign mem_MPORT_177_data = 20'h0;
  assign mem_MPORT_177_addr = 8'hb1;
  assign mem_MPORT_177_mask = 1'h1;
  assign mem_MPORT_177_en = reset;
  assign mem_MPORT_178_data = 20'h0;
  assign mem_MPORT_178_addr = 8'hb2;
  assign mem_MPORT_178_mask = 1'h1;
  assign mem_MPORT_178_en = reset;
  assign mem_MPORT_179_data = 20'h0;
  assign mem_MPORT_179_addr = 8'hb3;
  assign mem_MPORT_179_mask = 1'h1;
  assign mem_MPORT_179_en = reset;
  assign mem_MPORT_180_data = 20'h0;
  assign mem_MPORT_180_addr = 8'hb4;
  assign mem_MPORT_180_mask = 1'h1;
  assign mem_MPORT_180_en = reset;
  assign mem_MPORT_181_data = 20'h0;
  assign mem_MPORT_181_addr = 8'hb5;
  assign mem_MPORT_181_mask = 1'h1;
  assign mem_MPORT_181_en = reset;
  assign mem_MPORT_182_data = 20'h0;
  assign mem_MPORT_182_addr = 8'hb6;
  assign mem_MPORT_182_mask = 1'h1;
  assign mem_MPORT_182_en = reset;
  assign mem_MPORT_183_data = 20'h0;
  assign mem_MPORT_183_addr = 8'hb7;
  assign mem_MPORT_183_mask = 1'h1;
  assign mem_MPORT_183_en = reset;
  assign mem_MPORT_184_data = 20'h0;
  assign mem_MPORT_184_addr = 8'hb8;
  assign mem_MPORT_184_mask = 1'h1;
  assign mem_MPORT_184_en = reset;
  assign mem_MPORT_185_data = 20'h0;
  assign mem_MPORT_185_addr = 8'hb9;
  assign mem_MPORT_185_mask = 1'h1;
  assign mem_MPORT_185_en = reset;
  assign mem_MPORT_186_data = 20'h0;
  assign mem_MPORT_186_addr = 8'hba;
  assign mem_MPORT_186_mask = 1'h1;
  assign mem_MPORT_186_en = reset;
  assign mem_MPORT_187_data = 20'h0;
  assign mem_MPORT_187_addr = 8'hbb;
  assign mem_MPORT_187_mask = 1'h1;
  assign mem_MPORT_187_en = reset;
  assign mem_MPORT_188_data = 20'h0;
  assign mem_MPORT_188_addr = 8'hbc;
  assign mem_MPORT_188_mask = 1'h1;
  assign mem_MPORT_188_en = reset;
  assign mem_MPORT_189_data = 20'h0;
  assign mem_MPORT_189_addr = 8'hbd;
  assign mem_MPORT_189_mask = 1'h1;
  assign mem_MPORT_189_en = reset;
  assign mem_MPORT_190_data = 20'h0;
  assign mem_MPORT_190_addr = 8'hbe;
  assign mem_MPORT_190_mask = 1'h1;
  assign mem_MPORT_190_en = reset;
  assign mem_MPORT_191_data = 20'h0;
  assign mem_MPORT_191_addr = 8'hbf;
  assign mem_MPORT_191_mask = 1'h1;
  assign mem_MPORT_191_en = reset;
  assign mem_MPORT_192_data = 20'h0;
  assign mem_MPORT_192_addr = 8'hc0;
  assign mem_MPORT_192_mask = 1'h1;
  assign mem_MPORT_192_en = reset;
  assign mem_MPORT_193_data = 20'h0;
  assign mem_MPORT_193_addr = 8'hc1;
  assign mem_MPORT_193_mask = 1'h1;
  assign mem_MPORT_193_en = reset;
  assign mem_MPORT_194_data = 20'h0;
  assign mem_MPORT_194_addr = 8'hc2;
  assign mem_MPORT_194_mask = 1'h1;
  assign mem_MPORT_194_en = reset;
  assign mem_MPORT_195_data = 20'h0;
  assign mem_MPORT_195_addr = 8'hc3;
  assign mem_MPORT_195_mask = 1'h1;
  assign mem_MPORT_195_en = reset;
  assign mem_MPORT_196_data = 20'h0;
  assign mem_MPORT_196_addr = 8'hc4;
  assign mem_MPORT_196_mask = 1'h1;
  assign mem_MPORT_196_en = reset;
  assign mem_MPORT_197_data = 20'h0;
  assign mem_MPORT_197_addr = 8'hc5;
  assign mem_MPORT_197_mask = 1'h1;
  assign mem_MPORT_197_en = reset;
  assign mem_MPORT_198_data = 20'h0;
  assign mem_MPORT_198_addr = 8'hc6;
  assign mem_MPORT_198_mask = 1'h1;
  assign mem_MPORT_198_en = reset;
  assign mem_MPORT_199_data = 20'h0;
  assign mem_MPORT_199_addr = 8'hc7;
  assign mem_MPORT_199_mask = 1'h1;
  assign mem_MPORT_199_en = reset;
  assign mem_MPORT_200_data = 20'h0;
  assign mem_MPORT_200_addr = 8'hc8;
  assign mem_MPORT_200_mask = 1'h1;
  assign mem_MPORT_200_en = reset;
  assign mem_MPORT_201_data = 20'h0;
  assign mem_MPORT_201_addr = 8'hc9;
  assign mem_MPORT_201_mask = 1'h1;
  assign mem_MPORT_201_en = reset;
  assign mem_MPORT_202_data = 20'h0;
  assign mem_MPORT_202_addr = 8'hca;
  assign mem_MPORT_202_mask = 1'h1;
  assign mem_MPORT_202_en = reset;
  assign mem_MPORT_203_data = 20'h0;
  assign mem_MPORT_203_addr = 8'hcb;
  assign mem_MPORT_203_mask = 1'h1;
  assign mem_MPORT_203_en = reset;
  assign mem_MPORT_204_data = 20'h0;
  assign mem_MPORT_204_addr = 8'hcc;
  assign mem_MPORT_204_mask = 1'h1;
  assign mem_MPORT_204_en = reset;
  assign mem_MPORT_205_data = 20'h0;
  assign mem_MPORT_205_addr = 8'hcd;
  assign mem_MPORT_205_mask = 1'h1;
  assign mem_MPORT_205_en = reset;
  assign mem_MPORT_206_data = 20'h0;
  assign mem_MPORT_206_addr = 8'hce;
  assign mem_MPORT_206_mask = 1'h1;
  assign mem_MPORT_206_en = reset;
  assign mem_MPORT_207_data = 20'h0;
  assign mem_MPORT_207_addr = 8'hcf;
  assign mem_MPORT_207_mask = 1'h1;
  assign mem_MPORT_207_en = reset;
  assign mem_MPORT_208_data = 20'h0;
  assign mem_MPORT_208_addr = 8'hd0;
  assign mem_MPORT_208_mask = 1'h1;
  assign mem_MPORT_208_en = reset;
  assign mem_MPORT_209_data = 20'h0;
  assign mem_MPORT_209_addr = 8'hd1;
  assign mem_MPORT_209_mask = 1'h1;
  assign mem_MPORT_209_en = reset;
  assign mem_MPORT_210_data = 20'h0;
  assign mem_MPORT_210_addr = 8'hd2;
  assign mem_MPORT_210_mask = 1'h1;
  assign mem_MPORT_210_en = reset;
  assign mem_MPORT_211_data = 20'h0;
  assign mem_MPORT_211_addr = 8'hd3;
  assign mem_MPORT_211_mask = 1'h1;
  assign mem_MPORT_211_en = reset;
  assign mem_MPORT_212_data = 20'h0;
  assign mem_MPORT_212_addr = 8'hd4;
  assign mem_MPORT_212_mask = 1'h1;
  assign mem_MPORT_212_en = reset;
  assign mem_MPORT_213_data = 20'h0;
  assign mem_MPORT_213_addr = 8'hd5;
  assign mem_MPORT_213_mask = 1'h1;
  assign mem_MPORT_213_en = reset;
  assign mem_MPORT_214_data = 20'h0;
  assign mem_MPORT_214_addr = 8'hd6;
  assign mem_MPORT_214_mask = 1'h1;
  assign mem_MPORT_214_en = reset;
  assign mem_MPORT_215_data = 20'h0;
  assign mem_MPORT_215_addr = 8'hd7;
  assign mem_MPORT_215_mask = 1'h1;
  assign mem_MPORT_215_en = reset;
  assign mem_MPORT_216_data = 20'h0;
  assign mem_MPORT_216_addr = 8'hd8;
  assign mem_MPORT_216_mask = 1'h1;
  assign mem_MPORT_216_en = reset;
  assign mem_MPORT_217_data = 20'h0;
  assign mem_MPORT_217_addr = 8'hd9;
  assign mem_MPORT_217_mask = 1'h1;
  assign mem_MPORT_217_en = reset;
  assign mem_MPORT_218_data = 20'h0;
  assign mem_MPORT_218_addr = 8'hda;
  assign mem_MPORT_218_mask = 1'h1;
  assign mem_MPORT_218_en = reset;
  assign mem_MPORT_219_data = 20'h0;
  assign mem_MPORT_219_addr = 8'hdb;
  assign mem_MPORT_219_mask = 1'h1;
  assign mem_MPORT_219_en = reset;
  assign mem_MPORT_220_data = 20'h0;
  assign mem_MPORT_220_addr = 8'hdc;
  assign mem_MPORT_220_mask = 1'h1;
  assign mem_MPORT_220_en = reset;
  assign mem_MPORT_221_data = 20'h0;
  assign mem_MPORT_221_addr = 8'hdd;
  assign mem_MPORT_221_mask = 1'h1;
  assign mem_MPORT_221_en = reset;
  assign mem_MPORT_222_data = 20'h0;
  assign mem_MPORT_222_addr = 8'hde;
  assign mem_MPORT_222_mask = 1'h1;
  assign mem_MPORT_222_en = reset;
  assign mem_MPORT_223_data = 20'h0;
  assign mem_MPORT_223_addr = 8'hdf;
  assign mem_MPORT_223_mask = 1'h1;
  assign mem_MPORT_223_en = reset;
  assign mem_MPORT_224_data = 20'h0;
  assign mem_MPORT_224_addr = 8'he0;
  assign mem_MPORT_224_mask = 1'h1;
  assign mem_MPORT_224_en = reset;
  assign mem_MPORT_225_data = 20'h0;
  assign mem_MPORT_225_addr = 8'he1;
  assign mem_MPORT_225_mask = 1'h1;
  assign mem_MPORT_225_en = reset;
  assign mem_MPORT_226_data = 20'h0;
  assign mem_MPORT_226_addr = 8'he2;
  assign mem_MPORT_226_mask = 1'h1;
  assign mem_MPORT_226_en = reset;
  assign mem_MPORT_227_data = 20'h0;
  assign mem_MPORT_227_addr = 8'he3;
  assign mem_MPORT_227_mask = 1'h1;
  assign mem_MPORT_227_en = reset;
  assign mem_MPORT_228_data = 20'h0;
  assign mem_MPORT_228_addr = 8'he4;
  assign mem_MPORT_228_mask = 1'h1;
  assign mem_MPORT_228_en = reset;
  assign mem_MPORT_229_data = 20'h0;
  assign mem_MPORT_229_addr = 8'he5;
  assign mem_MPORT_229_mask = 1'h1;
  assign mem_MPORT_229_en = reset;
  assign mem_MPORT_230_data = 20'h0;
  assign mem_MPORT_230_addr = 8'he6;
  assign mem_MPORT_230_mask = 1'h1;
  assign mem_MPORT_230_en = reset;
  assign mem_MPORT_231_data = 20'h0;
  assign mem_MPORT_231_addr = 8'he7;
  assign mem_MPORT_231_mask = 1'h1;
  assign mem_MPORT_231_en = reset;
  assign mem_MPORT_232_data = 20'h0;
  assign mem_MPORT_232_addr = 8'he8;
  assign mem_MPORT_232_mask = 1'h1;
  assign mem_MPORT_232_en = reset;
  assign mem_MPORT_233_data = 20'h0;
  assign mem_MPORT_233_addr = 8'he9;
  assign mem_MPORT_233_mask = 1'h1;
  assign mem_MPORT_233_en = reset;
  assign mem_MPORT_234_data = 20'h0;
  assign mem_MPORT_234_addr = 8'hea;
  assign mem_MPORT_234_mask = 1'h1;
  assign mem_MPORT_234_en = reset;
  assign mem_MPORT_235_data = 20'h0;
  assign mem_MPORT_235_addr = 8'heb;
  assign mem_MPORT_235_mask = 1'h1;
  assign mem_MPORT_235_en = reset;
  assign mem_MPORT_236_data = 20'h0;
  assign mem_MPORT_236_addr = 8'hec;
  assign mem_MPORT_236_mask = 1'h1;
  assign mem_MPORT_236_en = reset;
  assign mem_MPORT_237_data = 20'h0;
  assign mem_MPORT_237_addr = 8'hed;
  assign mem_MPORT_237_mask = 1'h1;
  assign mem_MPORT_237_en = reset;
  assign mem_MPORT_238_data = 20'h0;
  assign mem_MPORT_238_addr = 8'hee;
  assign mem_MPORT_238_mask = 1'h1;
  assign mem_MPORT_238_en = reset;
  assign mem_MPORT_239_data = 20'h0;
  assign mem_MPORT_239_addr = 8'hef;
  assign mem_MPORT_239_mask = 1'h1;
  assign mem_MPORT_239_en = reset;
  assign mem_MPORT_240_data = 20'h0;
  assign mem_MPORT_240_addr = 8'hf0;
  assign mem_MPORT_240_mask = 1'h1;
  assign mem_MPORT_240_en = reset;
  assign mem_MPORT_241_data = 20'h0;
  assign mem_MPORT_241_addr = 8'hf1;
  assign mem_MPORT_241_mask = 1'h1;
  assign mem_MPORT_241_en = reset;
  assign mem_MPORT_242_data = 20'h0;
  assign mem_MPORT_242_addr = 8'hf2;
  assign mem_MPORT_242_mask = 1'h1;
  assign mem_MPORT_242_en = reset;
  assign mem_MPORT_243_data = 20'h0;
  assign mem_MPORT_243_addr = 8'hf3;
  assign mem_MPORT_243_mask = 1'h1;
  assign mem_MPORT_243_en = reset;
  assign mem_MPORT_244_data = 20'h0;
  assign mem_MPORT_244_addr = 8'hf4;
  assign mem_MPORT_244_mask = 1'h1;
  assign mem_MPORT_244_en = reset;
  assign mem_MPORT_245_data = 20'h0;
  assign mem_MPORT_245_addr = 8'hf5;
  assign mem_MPORT_245_mask = 1'h1;
  assign mem_MPORT_245_en = reset;
  assign mem_MPORT_246_data = 20'h0;
  assign mem_MPORT_246_addr = 8'hf6;
  assign mem_MPORT_246_mask = 1'h1;
  assign mem_MPORT_246_en = reset;
  assign mem_MPORT_247_data = 20'h0;
  assign mem_MPORT_247_addr = 8'hf7;
  assign mem_MPORT_247_mask = 1'h1;
  assign mem_MPORT_247_en = reset;
  assign mem_MPORT_248_data = 20'h0;
  assign mem_MPORT_248_addr = 8'hf8;
  assign mem_MPORT_248_mask = 1'h1;
  assign mem_MPORT_248_en = reset;
  assign mem_MPORT_249_data = 20'h0;
  assign mem_MPORT_249_addr = 8'hf9;
  assign mem_MPORT_249_mask = 1'h1;
  assign mem_MPORT_249_en = reset;
  assign mem_MPORT_250_data = 20'h0;
  assign mem_MPORT_250_addr = 8'hfa;
  assign mem_MPORT_250_mask = 1'h1;
  assign mem_MPORT_250_en = reset;
  assign mem_MPORT_251_data = 20'h0;
  assign mem_MPORT_251_addr = 8'hfb;
  assign mem_MPORT_251_mask = 1'h1;
  assign mem_MPORT_251_en = reset;
  assign mem_MPORT_252_data = 20'h0;
  assign mem_MPORT_252_addr = 8'hfc;
  assign mem_MPORT_252_mask = 1'h1;
  assign mem_MPORT_252_en = reset;
  assign mem_MPORT_253_data = 20'h0;
  assign mem_MPORT_253_addr = 8'hfd;
  assign mem_MPORT_253_mask = 1'h1;
  assign mem_MPORT_253_en = reset;
  assign mem_MPORT_254_data = 20'h0;
  assign mem_MPORT_254_addr = 8'hfe;
  assign mem_MPORT_254_mask = 1'h1;
  assign mem_MPORT_254_en = reset;
  assign mem_MPORT_255_data = 20'h0;
  assign mem_MPORT_255_addr = 8'hff;
  assign mem_MPORT_255_mask = 1'h1;
  assign mem_MPORT_255_en = reset;
  assign mem_MPORT_256_data = io_w_data;
  assign mem_MPORT_256_addr = io_w_addr;
  assign mem_MPORT_256_mask = 1'h1;
  assign mem_MPORT_256_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_129_en & mem_MPORT_129_mask) begin
      mem[mem_MPORT_129_addr] <= mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_130_en & mem_MPORT_130_mask) begin
      mem[mem_MPORT_130_addr] <= mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_131_en & mem_MPORT_131_mask) begin
      mem[mem_MPORT_131_addr] <= mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_132_en & mem_MPORT_132_mask) begin
      mem[mem_MPORT_132_addr] <= mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_133_en & mem_MPORT_133_mask) begin
      mem[mem_MPORT_133_addr] <= mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_134_en & mem_MPORT_134_mask) begin
      mem[mem_MPORT_134_addr] <= mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_135_en & mem_MPORT_135_mask) begin
      mem[mem_MPORT_135_addr] <= mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_136_en & mem_MPORT_136_mask) begin
      mem[mem_MPORT_136_addr] <= mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_137_en & mem_MPORT_137_mask) begin
      mem[mem_MPORT_137_addr] <= mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_138_en & mem_MPORT_138_mask) begin
      mem[mem_MPORT_138_addr] <= mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_139_en & mem_MPORT_139_mask) begin
      mem[mem_MPORT_139_addr] <= mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_140_en & mem_MPORT_140_mask) begin
      mem[mem_MPORT_140_addr] <= mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_141_en & mem_MPORT_141_mask) begin
      mem[mem_MPORT_141_addr] <= mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_142_en & mem_MPORT_142_mask) begin
      mem[mem_MPORT_142_addr] <= mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_143_en & mem_MPORT_143_mask) begin
      mem[mem_MPORT_143_addr] <= mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_144_en & mem_MPORT_144_mask) begin
      mem[mem_MPORT_144_addr] <= mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_145_en & mem_MPORT_145_mask) begin
      mem[mem_MPORT_145_addr] <= mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_146_en & mem_MPORT_146_mask) begin
      mem[mem_MPORT_146_addr] <= mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_147_en & mem_MPORT_147_mask) begin
      mem[mem_MPORT_147_addr] <= mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_148_en & mem_MPORT_148_mask) begin
      mem[mem_MPORT_148_addr] <= mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_149_en & mem_MPORT_149_mask) begin
      mem[mem_MPORT_149_addr] <= mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_150_en & mem_MPORT_150_mask) begin
      mem[mem_MPORT_150_addr] <= mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_151_en & mem_MPORT_151_mask) begin
      mem[mem_MPORT_151_addr] <= mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_152_en & mem_MPORT_152_mask) begin
      mem[mem_MPORT_152_addr] <= mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_153_en & mem_MPORT_153_mask) begin
      mem[mem_MPORT_153_addr] <= mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_154_en & mem_MPORT_154_mask) begin
      mem[mem_MPORT_154_addr] <= mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_155_en & mem_MPORT_155_mask) begin
      mem[mem_MPORT_155_addr] <= mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_156_en & mem_MPORT_156_mask) begin
      mem[mem_MPORT_156_addr] <= mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_157_en & mem_MPORT_157_mask) begin
      mem[mem_MPORT_157_addr] <= mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_158_en & mem_MPORT_158_mask) begin
      mem[mem_MPORT_158_addr] <= mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_159_en & mem_MPORT_159_mask) begin
      mem[mem_MPORT_159_addr] <= mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_160_en & mem_MPORT_160_mask) begin
      mem[mem_MPORT_160_addr] <= mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_161_en & mem_MPORT_161_mask) begin
      mem[mem_MPORT_161_addr] <= mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_162_en & mem_MPORT_162_mask) begin
      mem[mem_MPORT_162_addr] <= mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_163_en & mem_MPORT_163_mask) begin
      mem[mem_MPORT_163_addr] <= mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_164_en & mem_MPORT_164_mask) begin
      mem[mem_MPORT_164_addr] <= mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_165_en & mem_MPORT_165_mask) begin
      mem[mem_MPORT_165_addr] <= mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_166_en & mem_MPORT_166_mask) begin
      mem[mem_MPORT_166_addr] <= mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_167_en & mem_MPORT_167_mask) begin
      mem[mem_MPORT_167_addr] <= mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_168_en & mem_MPORT_168_mask) begin
      mem[mem_MPORT_168_addr] <= mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_169_en & mem_MPORT_169_mask) begin
      mem[mem_MPORT_169_addr] <= mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_170_en & mem_MPORT_170_mask) begin
      mem[mem_MPORT_170_addr] <= mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_171_en & mem_MPORT_171_mask) begin
      mem[mem_MPORT_171_addr] <= mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_172_en & mem_MPORT_172_mask) begin
      mem[mem_MPORT_172_addr] <= mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_173_en & mem_MPORT_173_mask) begin
      mem[mem_MPORT_173_addr] <= mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_174_en & mem_MPORT_174_mask) begin
      mem[mem_MPORT_174_addr] <= mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_175_en & mem_MPORT_175_mask) begin
      mem[mem_MPORT_175_addr] <= mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_176_en & mem_MPORT_176_mask) begin
      mem[mem_MPORT_176_addr] <= mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_177_en & mem_MPORT_177_mask) begin
      mem[mem_MPORT_177_addr] <= mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_178_en & mem_MPORT_178_mask) begin
      mem[mem_MPORT_178_addr] <= mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_179_en & mem_MPORT_179_mask) begin
      mem[mem_MPORT_179_addr] <= mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_180_en & mem_MPORT_180_mask) begin
      mem[mem_MPORT_180_addr] <= mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_181_en & mem_MPORT_181_mask) begin
      mem[mem_MPORT_181_addr] <= mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_182_en & mem_MPORT_182_mask) begin
      mem[mem_MPORT_182_addr] <= mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_183_en & mem_MPORT_183_mask) begin
      mem[mem_MPORT_183_addr] <= mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_184_en & mem_MPORT_184_mask) begin
      mem[mem_MPORT_184_addr] <= mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_185_en & mem_MPORT_185_mask) begin
      mem[mem_MPORT_185_addr] <= mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_186_en & mem_MPORT_186_mask) begin
      mem[mem_MPORT_186_addr] <= mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_187_en & mem_MPORT_187_mask) begin
      mem[mem_MPORT_187_addr] <= mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_188_en & mem_MPORT_188_mask) begin
      mem[mem_MPORT_188_addr] <= mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_189_en & mem_MPORT_189_mask) begin
      mem[mem_MPORT_189_addr] <= mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_190_en & mem_MPORT_190_mask) begin
      mem[mem_MPORT_190_addr] <= mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_191_en & mem_MPORT_191_mask) begin
      mem[mem_MPORT_191_addr] <= mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_192_en & mem_MPORT_192_mask) begin
      mem[mem_MPORT_192_addr] <= mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_193_en & mem_MPORT_193_mask) begin
      mem[mem_MPORT_193_addr] <= mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_194_en & mem_MPORT_194_mask) begin
      mem[mem_MPORT_194_addr] <= mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_195_en & mem_MPORT_195_mask) begin
      mem[mem_MPORT_195_addr] <= mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_196_en & mem_MPORT_196_mask) begin
      mem[mem_MPORT_196_addr] <= mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_197_en & mem_MPORT_197_mask) begin
      mem[mem_MPORT_197_addr] <= mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_198_en & mem_MPORT_198_mask) begin
      mem[mem_MPORT_198_addr] <= mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_199_en & mem_MPORT_199_mask) begin
      mem[mem_MPORT_199_addr] <= mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_200_en & mem_MPORT_200_mask) begin
      mem[mem_MPORT_200_addr] <= mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_201_en & mem_MPORT_201_mask) begin
      mem[mem_MPORT_201_addr] <= mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_202_en & mem_MPORT_202_mask) begin
      mem[mem_MPORT_202_addr] <= mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_203_en & mem_MPORT_203_mask) begin
      mem[mem_MPORT_203_addr] <= mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_204_en & mem_MPORT_204_mask) begin
      mem[mem_MPORT_204_addr] <= mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_205_en & mem_MPORT_205_mask) begin
      mem[mem_MPORT_205_addr] <= mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_206_en & mem_MPORT_206_mask) begin
      mem[mem_MPORT_206_addr] <= mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_207_en & mem_MPORT_207_mask) begin
      mem[mem_MPORT_207_addr] <= mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_208_en & mem_MPORT_208_mask) begin
      mem[mem_MPORT_208_addr] <= mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_209_en & mem_MPORT_209_mask) begin
      mem[mem_MPORT_209_addr] <= mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_210_en & mem_MPORT_210_mask) begin
      mem[mem_MPORT_210_addr] <= mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_211_en & mem_MPORT_211_mask) begin
      mem[mem_MPORT_211_addr] <= mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_212_en & mem_MPORT_212_mask) begin
      mem[mem_MPORT_212_addr] <= mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_213_en & mem_MPORT_213_mask) begin
      mem[mem_MPORT_213_addr] <= mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_214_en & mem_MPORT_214_mask) begin
      mem[mem_MPORT_214_addr] <= mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_215_en & mem_MPORT_215_mask) begin
      mem[mem_MPORT_215_addr] <= mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_216_en & mem_MPORT_216_mask) begin
      mem[mem_MPORT_216_addr] <= mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_217_en & mem_MPORT_217_mask) begin
      mem[mem_MPORT_217_addr] <= mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_218_en & mem_MPORT_218_mask) begin
      mem[mem_MPORT_218_addr] <= mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_219_en & mem_MPORT_219_mask) begin
      mem[mem_MPORT_219_addr] <= mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_220_en & mem_MPORT_220_mask) begin
      mem[mem_MPORT_220_addr] <= mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_221_en & mem_MPORT_221_mask) begin
      mem[mem_MPORT_221_addr] <= mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_222_en & mem_MPORT_222_mask) begin
      mem[mem_MPORT_222_addr] <= mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_223_en & mem_MPORT_223_mask) begin
      mem[mem_MPORT_223_addr] <= mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_224_en & mem_MPORT_224_mask) begin
      mem[mem_MPORT_224_addr] <= mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_225_en & mem_MPORT_225_mask) begin
      mem[mem_MPORT_225_addr] <= mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_226_en & mem_MPORT_226_mask) begin
      mem[mem_MPORT_226_addr] <= mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_227_en & mem_MPORT_227_mask) begin
      mem[mem_MPORT_227_addr] <= mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_228_en & mem_MPORT_228_mask) begin
      mem[mem_MPORT_228_addr] <= mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_229_en & mem_MPORT_229_mask) begin
      mem[mem_MPORT_229_addr] <= mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_230_en & mem_MPORT_230_mask) begin
      mem[mem_MPORT_230_addr] <= mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_231_en & mem_MPORT_231_mask) begin
      mem[mem_MPORT_231_addr] <= mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_232_en & mem_MPORT_232_mask) begin
      mem[mem_MPORT_232_addr] <= mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_233_en & mem_MPORT_233_mask) begin
      mem[mem_MPORT_233_addr] <= mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_234_en & mem_MPORT_234_mask) begin
      mem[mem_MPORT_234_addr] <= mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_235_en & mem_MPORT_235_mask) begin
      mem[mem_MPORT_235_addr] <= mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_236_en & mem_MPORT_236_mask) begin
      mem[mem_MPORT_236_addr] <= mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_237_en & mem_MPORT_237_mask) begin
      mem[mem_MPORT_237_addr] <= mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_238_en & mem_MPORT_238_mask) begin
      mem[mem_MPORT_238_addr] <= mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_239_en & mem_MPORT_239_mask) begin
      mem[mem_MPORT_239_addr] <= mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_240_en & mem_MPORT_240_mask) begin
      mem[mem_MPORT_240_addr] <= mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_241_en & mem_MPORT_241_mask) begin
      mem[mem_MPORT_241_addr] <= mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_242_en & mem_MPORT_242_mask) begin
      mem[mem_MPORT_242_addr] <= mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_243_en & mem_MPORT_243_mask) begin
      mem[mem_MPORT_243_addr] <= mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_244_en & mem_MPORT_244_mask) begin
      mem[mem_MPORT_244_addr] <= mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_245_en & mem_MPORT_245_mask) begin
      mem[mem_MPORT_245_addr] <= mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_246_en & mem_MPORT_246_mask) begin
      mem[mem_MPORT_246_addr] <= mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_247_en & mem_MPORT_247_mask) begin
      mem[mem_MPORT_247_addr] <= mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_248_en & mem_MPORT_248_mask) begin
      mem[mem_MPORT_248_addr] <= mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_249_en & mem_MPORT_249_mask) begin
      mem[mem_MPORT_249_addr] <= mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_250_en & mem_MPORT_250_mask) begin
      mem[mem_MPORT_250_addr] <= mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_251_en & mem_MPORT_251_mask) begin
      mem[mem_MPORT_251_addr] <= mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_252_en & mem_MPORT_252_mask) begin
      mem[mem_MPORT_252_addr] <= mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_253_en & mem_MPORT_253_mask) begin
      mem[mem_MPORT_253_addr] <= mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_254_en & mem_MPORT_254_mask) begin
      mem[mem_MPORT_254_addr] <= mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_255_en & mem_MPORT_255_mask) begin
      mem[mem_MPORT_255_addr] <= mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_256_en & mem_MPORT_256_mask) begin
      mem[mem_MPORT_256_addr] <= mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _RAND_0[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_18(
  input         clock,
  input         reset,
  input  [7:0]  io_r_addr,
  output [19:0] io_r_data_0,
  output [19:0] io_r_data_1,
  output [19:0] io_r_data_2,
  output [19:0] io_r_data_3,
  output [19:0] io_r_data_4,
  output [19:0] io_r_data_5,
  output [19:0] io_r_data_6,
  output [19:0] io_r_data_7,
  input         io_w_en,
  input  [7:0]  io_w_addr,
  input  [19:0] io_w_data_0,
  input  [19:0] io_w_data_1,
  input  [19:0] io_w_data_2,
  input  [19:0] io_w_data_3,
  input  [19:0] io_w_data_4,
  input  [19:0] io_w_data_5,
  input  [19:0] io_w_data_6,
  input  [19:0] io_w_data_7,
  input  [7:0]  io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_clock; // @[SRAM_1.scala 201:38]
  wire  brams_4_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_4_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_4_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_4_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_4_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_clock; // @[SRAM_1.scala 201:38]
  wire  brams_5_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_5_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_5_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_5_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_5_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_clock; // @[SRAM_1.scala 201:38]
  wire  brams_6_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_6_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_6_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_6_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_6_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_clock; // @[SRAM_1.scala 201:38]
  wire  brams_7_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_7_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_7_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_7_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [19:0] brams_7_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P_112 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P_112 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P_112 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P_112 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  BankRAM_2P_112 brams_4 ( // @[SRAM_1.scala 201:38]
    .clock(brams_4_clock),
    .reset(brams_4_reset),
    .io_r_addr(brams_4_io_r_addr),
    .io_r_data(brams_4_io_r_data),
    .io_w_en(brams_4_io_w_en),
    .io_w_addr(brams_4_io_w_addr),
    .io_w_data(brams_4_io_w_data)
  );
  BankRAM_2P_112 brams_5 ( // @[SRAM_1.scala 201:38]
    .clock(brams_5_clock),
    .reset(brams_5_reset),
    .io_r_addr(brams_5_io_r_addr),
    .io_r_data(brams_5_io_r_data),
    .io_w_en(brams_5_io_w_en),
    .io_w_addr(brams_5_io_w_addr),
    .io_w_data(brams_5_io_w_data)
  );
  BankRAM_2P_112 brams_6 ( // @[SRAM_1.scala 201:38]
    .clock(brams_6_clock),
    .reset(brams_6_reset),
    .io_r_addr(brams_6_io_r_addr),
    .io_r_data(brams_6_io_r_data),
    .io_w_en(brams_6_io_w_en),
    .io_w_addr(brams_6_io_w_addr),
    .io_w_data(brams_6_io_w_data)
  );
  BankRAM_2P_112 brams_7 ( // @[SRAM_1.scala 201:38]
    .clock(brams_7_clock),
    .reset(brams_7_reset),
    .io_r_addr(brams_7_io_r_addr),
    .io_r_data(brams_7_io_r_data),
    .io_w_en(brams_7_io_w_en),
    .io_w_addr(brams_7_io_w_addr),
    .io_w_data(brams_7_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_4 = brams_4_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_5 = brams_5_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_6 = brams_6_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_7 = brams_7_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
  assign brams_4_clock = clock;
  assign brams_4_reset = reset;
  assign brams_4_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_4_io_w_en = io_w_en & io_w_maskOH[4]; // @[SRAM_1.scala 208:37]
  assign brams_4_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_4_io_w_data = io_w_data_4; // @[SRAM_1.scala 210:28]
  assign brams_5_clock = clock;
  assign brams_5_reset = reset;
  assign brams_5_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_5_io_w_en = io_w_en & io_w_maskOH[5]; // @[SRAM_1.scala 208:37]
  assign brams_5_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_5_io_w_data = io_w_data_5; // @[SRAM_1.scala 210:28]
  assign brams_6_clock = clock;
  assign brams_6_reset = reset;
  assign brams_6_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_6_io_w_en = io_w_en & io_w_maskOH[6]; // @[SRAM_1.scala 208:37]
  assign brams_6_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_6_io_w_data = io_w_data_6; // @[SRAM_1.scala 210:28]
  assign brams_7_clock = clock;
  assign brams_7_reset = reset;
  assign brams_7_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_7_io_w_en = io_w_en & io_w_maskOH[7]; // @[SRAM_1.scala 208:37]
  assign brams_7_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_7_io_w_data = io_w_data_7; // @[SRAM_1.scala 210:28]
endmodule
module BankRAM_2P_120(
  input        clock,
  input        reset,
  input  [7:0] io_r_addr,
  output [1:0] io_r_data,
  input        io_w_en,
  input  [7:0] io_w_addr,
  input  [1:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] mem [0:255]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_129_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_130_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_131_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_132_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_133_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_134_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_135_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_136_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_137_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_138_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_139_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_140_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_141_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_142_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_143_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_144_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_145_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_146_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_147_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_148_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_149_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_150_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_151_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_152_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_153_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_154_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_155_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_156_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_157_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_158_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_159_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_160_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_161_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_162_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_163_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_164_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_165_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_166_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_167_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_168_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_169_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_170_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_171_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_172_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_173_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_174_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_175_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_176_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_177_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_178_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_179_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_180_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_181_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_182_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_183_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_184_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_185_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_186_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_187_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_188_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_189_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_190_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_191_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_192_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_193_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_194_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_195_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_196_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_197_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_198_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_199_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_200_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_201_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_202_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_203_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_204_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_205_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_206_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_207_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_208_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_209_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_210_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_211_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_212_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_213_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_214_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_215_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_216_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_217_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_218_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_219_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_220_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_221_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_222_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_223_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_224_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_225_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_226_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_227_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_228_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_229_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_230_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_231_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_232_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_233_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_234_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_235_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_236_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_237_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_238_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_239_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_240_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_241_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_242_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_243_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_244_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_245_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_246_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_247_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_248_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_249_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_250_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_251_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_252_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_253_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_254_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_255_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
  wire [7:0] mem_MPORT_256_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [7:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 2'h0;
  assign mem_MPORT_addr = 8'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 2'h0;
  assign mem_MPORT_1_addr = 8'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 2'h0;
  assign mem_MPORT_2_addr = 8'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 2'h0;
  assign mem_MPORT_3_addr = 8'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 2'h0;
  assign mem_MPORT_4_addr = 8'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 2'h0;
  assign mem_MPORT_5_addr = 8'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 2'h0;
  assign mem_MPORT_6_addr = 8'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 2'h0;
  assign mem_MPORT_7_addr = 8'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 2'h0;
  assign mem_MPORT_8_addr = 8'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 2'h0;
  assign mem_MPORT_9_addr = 8'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 2'h0;
  assign mem_MPORT_10_addr = 8'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 2'h0;
  assign mem_MPORT_11_addr = 8'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 2'h0;
  assign mem_MPORT_12_addr = 8'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 2'h0;
  assign mem_MPORT_13_addr = 8'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 2'h0;
  assign mem_MPORT_14_addr = 8'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 2'h0;
  assign mem_MPORT_15_addr = 8'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 2'h0;
  assign mem_MPORT_16_addr = 8'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 2'h0;
  assign mem_MPORT_17_addr = 8'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 2'h0;
  assign mem_MPORT_18_addr = 8'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 2'h0;
  assign mem_MPORT_19_addr = 8'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 2'h0;
  assign mem_MPORT_20_addr = 8'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 2'h0;
  assign mem_MPORT_21_addr = 8'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 2'h0;
  assign mem_MPORT_22_addr = 8'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 2'h0;
  assign mem_MPORT_23_addr = 8'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 2'h0;
  assign mem_MPORT_24_addr = 8'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 2'h0;
  assign mem_MPORT_25_addr = 8'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 2'h0;
  assign mem_MPORT_26_addr = 8'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 2'h0;
  assign mem_MPORT_27_addr = 8'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 2'h0;
  assign mem_MPORT_28_addr = 8'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 2'h0;
  assign mem_MPORT_29_addr = 8'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 2'h0;
  assign mem_MPORT_30_addr = 8'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 2'h0;
  assign mem_MPORT_31_addr = 8'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 2'h0;
  assign mem_MPORT_32_addr = 8'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 2'h0;
  assign mem_MPORT_33_addr = 8'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 2'h0;
  assign mem_MPORT_34_addr = 8'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 2'h0;
  assign mem_MPORT_35_addr = 8'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 2'h0;
  assign mem_MPORT_36_addr = 8'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 2'h0;
  assign mem_MPORT_37_addr = 8'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 2'h0;
  assign mem_MPORT_38_addr = 8'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 2'h0;
  assign mem_MPORT_39_addr = 8'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 2'h0;
  assign mem_MPORT_40_addr = 8'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 2'h0;
  assign mem_MPORT_41_addr = 8'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 2'h0;
  assign mem_MPORT_42_addr = 8'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 2'h0;
  assign mem_MPORT_43_addr = 8'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 2'h0;
  assign mem_MPORT_44_addr = 8'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 2'h0;
  assign mem_MPORT_45_addr = 8'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 2'h0;
  assign mem_MPORT_46_addr = 8'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 2'h0;
  assign mem_MPORT_47_addr = 8'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 2'h0;
  assign mem_MPORT_48_addr = 8'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 2'h0;
  assign mem_MPORT_49_addr = 8'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 2'h0;
  assign mem_MPORT_50_addr = 8'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 2'h0;
  assign mem_MPORT_51_addr = 8'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 2'h0;
  assign mem_MPORT_52_addr = 8'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 2'h0;
  assign mem_MPORT_53_addr = 8'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 2'h0;
  assign mem_MPORT_54_addr = 8'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 2'h0;
  assign mem_MPORT_55_addr = 8'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 2'h0;
  assign mem_MPORT_56_addr = 8'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 2'h0;
  assign mem_MPORT_57_addr = 8'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 2'h0;
  assign mem_MPORT_58_addr = 8'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 2'h0;
  assign mem_MPORT_59_addr = 8'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 2'h0;
  assign mem_MPORT_60_addr = 8'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 2'h0;
  assign mem_MPORT_61_addr = 8'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 2'h0;
  assign mem_MPORT_62_addr = 8'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 2'h0;
  assign mem_MPORT_63_addr = 8'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 2'h0;
  assign mem_MPORT_64_addr = 8'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 2'h0;
  assign mem_MPORT_65_addr = 8'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 2'h0;
  assign mem_MPORT_66_addr = 8'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 2'h0;
  assign mem_MPORT_67_addr = 8'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 2'h0;
  assign mem_MPORT_68_addr = 8'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 2'h0;
  assign mem_MPORT_69_addr = 8'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 2'h0;
  assign mem_MPORT_70_addr = 8'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 2'h0;
  assign mem_MPORT_71_addr = 8'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 2'h0;
  assign mem_MPORT_72_addr = 8'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 2'h0;
  assign mem_MPORT_73_addr = 8'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 2'h0;
  assign mem_MPORT_74_addr = 8'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 2'h0;
  assign mem_MPORT_75_addr = 8'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 2'h0;
  assign mem_MPORT_76_addr = 8'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 2'h0;
  assign mem_MPORT_77_addr = 8'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 2'h0;
  assign mem_MPORT_78_addr = 8'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 2'h0;
  assign mem_MPORT_79_addr = 8'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 2'h0;
  assign mem_MPORT_80_addr = 8'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 2'h0;
  assign mem_MPORT_81_addr = 8'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 2'h0;
  assign mem_MPORT_82_addr = 8'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 2'h0;
  assign mem_MPORT_83_addr = 8'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 2'h0;
  assign mem_MPORT_84_addr = 8'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 2'h0;
  assign mem_MPORT_85_addr = 8'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 2'h0;
  assign mem_MPORT_86_addr = 8'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 2'h0;
  assign mem_MPORT_87_addr = 8'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 2'h0;
  assign mem_MPORT_88_addr = 8'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 2'h0;
  assign mem_MPORT_89_addr = 8'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 2'h0;
  assign mem_MPORT_90_addr = 8'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 2'h0;
  assign mem_MPORT_91_addr = 8'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 2'h0;
  assign mem_MPORT_92_addr = 8'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 2'h0;
  assign mem_MPORT_93_addr = 8'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 2'h0;
  assign mem_MPORT_94_addr = 8'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 2'h0;
  assign mem_MPORT_95_addr = 8'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 2'h0;
  assign mem_MPORT_96_addr = 8'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 2'h0;
  assign mem_MPORT_97_addr = 8'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 2'h0;
  assign mem_MPORT_98_addr = 8'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 2'h0;
  assign mem_MPORT_99_addr = 8'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 2'h0;
  assign mem_MPORT_100_addr = 8'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 2'h0;
  assign mem_MPORT_101_addr = 8'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 2'h0;
  assign mem_MPORT_102_addr = 8'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 2'h0;
  assign mem_MPORT_103_addr = 8'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 2'h0;
  assign mem_MPORT_104_addr = 8'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 2'h0;
  assign mem_MPORT_105_addr = 8'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 2'h0;
  assign mem_MPORT_106_addr = 8'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 2'h0;
  assign mem_MPORT_107_addr = 8'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 2'h0;
  assign mem_MPORT_108_addr = 8'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 2'h0;
  assign mem_MPORT_109_addr = 8'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 2'h0;
  assign mem_MPORT_110_addr = 8'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 2'h0;
  assign mem_MPORT_111_addr = 8'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 2'h0;
  assign mem_MPORT_112_addr = 8'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 2'h0;
  assign mem_MPORT_113_addr = 8'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 2'h0;
  assign mem_MPORT_114_addr = 8'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 2'h0;
  assign mem_MPORT_115_addr = 8'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 2'h0;
  assign mem_MPORT_116_addr = 8'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 2'h0;
  assign mem_MPORT_117_addr = 8'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 2'h0;
  assign mem_MPORT_118_addr = 8'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 2'h0;
  assign mem_MPORT_119_addr = 8'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 2'h0;
  assign mem_MPORT_120_addr = 8'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 2'h0;
  assign mem_MPORT_121_addr = 8'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 2'h0;
  assign mem_MPORT_122_addr = 8'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 2'h0;
  assign mem_MPORT_123_addr = 8'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 2'h0;
  assign mem_MPORT_124_addr = 8'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 2'h0;
  assign mem_MPORT_125_addr = 8'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 2'h0;
  assign mem_MPORT_126_addr = 8'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 2'h0;
  assign mem_MPORT_127_addr = 8'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 2'h0;
  assign mem_MPORT_128_addr = 8'h80;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = reset;
  assign mem_MPORT_129_data = 2'h0;
  assign mem_MPORT_129_addr = 8'h81;
  assign mem_MPORT_129_mask = 1'h1;
  assign mem_MPORT_129_en = reset;
  assign mem_MPORT_130_data = 2'h0;
  assign mem_MPORT_130_addr = 8'h82;
  assign mem_MPORT_130_mask = 1'h1;
  assign mem_MPORT_130_en = reset;
  assign mem_MPORT_131_data = 2'h0;
  assign mem_MPORT_131_addr = 8'h83;
  assign mem_MPORT_131_mask = 1'h1;
  assign mem_MPORT_131_en = reset;
  assign mem_MPORT_132_data = 2'h0;
  assign mem_MPORT_132_addr = 8'h84;
  assign mem_MPORT_132_mask = 1'h1;
  assign mem_MPORT_132_en = reset;
  assign mem_MPORT_133_data = 2'h0;
  assign mem_MPORT_133_addr = 8'h85;
  assign mem_MPORT_133_mask = 1'h1;
  assign mem_MPORT_133_en = reset;
  assign mem_MPORT_134_data = 2'h0;
  assign mem_MPORT_134_addr = 8'h86;
  assign mem_MPORT_134_mask = 1'h1;
  assign mem_MPORT_134_en = reset;
  assign mem_MPORT_135_data = 2'h0;
  assign mem_MPORT_135_addr = 8'h87;
  assign mem_MPORT_135_mask = 1'h1;
  assign mem_MPORT_135_en = reset;
  assign mem_MPORT_136_data = 2'h0;
  assign mem_MPORT_136_addr = 8'h88;
  assign mem_MPORT_136_mask = 1'h1;
  assign mem_MPORT_136_en = reset;
  assign mem_MPORT_137_data = 2'h0;
  assign mem_MPORT_137_addr = 8'h89;
  assign mem_MPORT_137_mask = 1'h1;
  assign mem_MPORT_137_en = reset;
  assign mem_MPORT_138_data = 2'h0;
  assign mem_MPORT_138_addr = 8'h8a;
  assign mem_MPORT_138_mask = 1'h1;
  assign mem_MPORT_138_en = reset;
  assign mem_MPORT_139_data = 2'h0;
  assign mem_MPORT_139_addr = 8'h8b;
  assign mem_MPORT_139_mask = 1'h1;
  assign mem_MPORT_139_en = reset;
  assign mem_MPORT_140_data = 2'h0;
  assign mem_MPORT_140_addr = 8'h8c;
  assign mem_MPORT_140_mask = 1'h1;
  assign mem_MPORT_140_en = reset;
  assign mem_MPORT_141_data = 2'h0;
  assign mem_MPORT_141_addr = 8'h8d;
  assign mem_MPORT_141_mask = 1'h1;
  assign mem_MPORT_141_en = reset;
  assign mem_MPORT_142_data = 2'h0;
  assign mem_MPORT_142_addr = 8'h8e;
  assign mem_MPORT_142_mask = 1'h1;
  assign mem_MPORT_142_en = reset;
  assign mem_MPORT_143_data = 2'h0;
  assign mem_MPORT_143_addr = 8'h8f;
  assign mem_MPORT_143_mask = 1'h1;
  assign mem_MPORT_143_en = reset;
  assign mem_MPORT_144_data = 2'h0;
  assign mem_MPORT_144_addr = 8'h90;
  assign mem_MPORT_144_mask = 1'h1;
  assign mem_MPORT_144_en = reset;
  assign mem_MPORT_145_data = 2'h0;
  assign mem_MPORT_145_addr = 8'h91;
  assign mem_MPORT_145_mask = 1'h1;
  assign mem_MPORT_145_en = reset;
  assign mem_MPORT_146_data = 2'h0;
  assign mem_MPORT_146_addr = 8'h92;
  assign mem_MPORT_146_mask = 1'h1;
  assign mem_MPORT_146_en = reset;
  assign mem_MPORT_147_data = 2'h0;
  assign mem_MPORT_147_addr = 8'h93;
  assign mem_MPORT_147_mask = 1'h1;
  assign mem_MPORT_147_en = reset;
  assign mem_MPORT_148_data = 2'h0;
  assign mem_MPORT_148_addr = 8'h94;
  assign mem_MPORT_148_mask = 1'h1;
  assign mem_MPORT_148_en = reset;
  assign mem_MPORT_149_data = 2'h0;
  assign mem_MPORT_149_addr = 8'h95;
  assign mem_MPORT_149_mask = 1'h1;
  assign mem_MPORT_149_en = reset;
  assign mem_MPORT_150_data = 2'h0;
  assign mem_MPORT_150_addr = 8'h96;
  assign mem_MPORT_150_mask = 1'h1;
  assign mem_MPORT_150_en = reset;
  assign mem_MPORT_151_data = 2'h0;
  assign mem_MPORT_151_addr = 8'h97;
  assign mem_MPORT_151_mask = 1'h1;
  assign mem_MPORT_151_en = reset;
  assign mem_MPORT_152_data = 2'h0;
  assign mem_MPORT_152_addr = 8'h98;
  assign mem_MPORT_152_mask = 1'h1;
  assign mem_MPORT_152_en = reset;
  assign mem_MPORT_153_data = 2'h0;
  assign mem_MPORT_153_addr = 8'h99;
  assign mem_MPORT_153_mask = 1'h1;
  assign mem_MPORT_153_en = reset;
  assign mem_MPORT_154_data = 2'h0;
  assign mem_MPORT_154_addr = 8'h9a;
  assign mem_MPORT_154_mask = 1'h1;
  assign mem_MPORT_154_en = reset;
  assign mem_MPORT_155_data = 2'h0;
  assign mem_MPORT_155_addr = 8'h9b;
  assign mem_MPORT_155_mask = 1'h1;
  assign mem_MPORT_155_en = reset;
  assign mem_MPORT_156_data = 2'h0;
  assign mem_MPORT_156_addr = 8'h9c;
  assign mem_MPORT_156_mask = 1'h1;
  assign mem_MPORT_156_en = reset;
  assign mem_MPORT_157_data = 2'h0;
  assign mem_MPORT_157_addr = 8'h9d;
  assign mem_MPORT_157_mask = 1'h1;
  assign mem_MPORT_157_en = reset;
  assign mem_MPORT_158_data = 2'h0;
  assign mem_MPORT_158_addr = 8'h9e;
  assign mem_MPORT_158_mask = 1'h1;
  assign mem_MPORT_158_en = reset;
  assign mem_MPORT_159_data = 2'h0;
  assign mem_MPORT_159_addr = 8'h9f;
  assign mem_MPORT_159_mask = 1'h1;
  assign mem_MPORT_159_en = reset;
  assign mem_MPORT_160_data = 2'h0;
  assign mem_MPORT_160_addr = 8'ha0;
  assign mem_MPORT_160_mask = 1'h1;
  assign mem_MPORT_160_en = reset;
  assign mem_MPORT_161_data = 2'h0;
  assign mem_MPORT_161_addr = 8'ha1;
  assign mem_MPORT_161_mask = 1'h1;
  assign mem_MPORT_161_en = reset;
  assign mem_MPORT_162_data = 2'h0;
  assign mem_MPORT_162_addr = 8'ha2;
  assign mem_MPORT_162_mask = 1'h1;
  assign mem_MPORT_162_en = reset;
  assign mem_MPORT_163_data = 2'h0;
  assign mem_MPORT_163_addr = 8'ha3;
  assign mem_MPORT_163_mask = 1'h1;
  assign mem_MPORT_163_en = reset;
  assign mem_MPORT_164_data = 2'h0;
  assign mem_MPORT_164_addr = 8'ha4;
  assign mem_MPORT_164_mask = 1'h1;
  assign mem_MPORT_164_en = reset;
  assign mem_MPORT_165_data = 2'h0;
  assign mem_MPORT_165_addr = 8'ha5;
  assign mem_MPORT_165_mask = 1'h1;
  assign mem_MPORT_165_en = reset;
  assign mem_MPORT_166_data = 2'h0;
  assign mem_MPORT_166_addr = 8'ha6;
  assign mem_MPORT_166_mask = 1'h1;
  assign mem_MPORT_166_en = reset;
  assign mem_MPORT_167_data = 2'h0;
  assign mem_MPORT_167_addr = 8'ha7;
  assign mem_MPORT_167_mask = 1'h1;
  assign mem_MPORT_167_en = reset;
  assign mem_MPORT_168_data = 2'h0;
  assign mem_MPORT_168_addr = 8'ha8;
  assign mem_MPORT_168_mask = 1'h1;
  assign mem_MPORT_168_en = reset;
  assign mem_MPORT_169_data = 2'h0;
  assign mem_MPORT_169_addr = 8'ha9;
  assign mem_MPORT_169_mask = 1'h1;
  assign mem_MPORT_169_en = reset;
  assign mem_MPORT_170_data = 2'h0;
  assign mem_MPORT_170_addr = 8'haa;
  assign mem_MPORT_170_mask = 1'h1;
  assign mem_MPORT_170_en = reset;
  assign mem_MPORT_171_data = 2'h0;
  assign mem_MPORT_171_addr = 8'hab;
  assign mem_MPORT_171_mask = 1'h1;
  assign mem_MPORT_171_en = reset;
  assign mem_MPORT_172_data = 2'h0;
  assign mem_MPORT_172_addr = 8'hac;
  assign mem_MPORT_172_mask = 1'h1;
  assign mem_MPORT_172_en = reset;
  assign mem_MPORT_173_data = 2'h0;
  assign mem_MPORT_173_addr = 8'had;
  assign mem_MPORT_173_mask = 1'h1;
  assign mem_MPORT_173_en = reset;
  assign mem_MPORT_174_data = 2'h0;
  assign mem_MPORT_174_addr = 8'hae;
  assign mem_MPORT_174_mask = 1'h1;
  assign mem_MPORT_174_en = reset;
  assign mem_MPORT_175_data = 2'h0;
  assign mem_MPORT_175_addr = 8'haf;
  assign mem_MPORT_175_mask = 1'h1;
  assign mem_MPORT_175_en = reset;
  assign mem_MPORT_176_data = 2'h0;
  assign mem_MPORT_176_addr = 8'hb0;
  assign mem_MPORT_176_mask = 1'h1;
  assign mem_MPORT_176_en = reset;
  assign mem_MPORT_177_data = 2'h0;
  assign mem_MPORT_177_addr = 8'hb1;
  assign mem_MPORT_177_mask = 1'h1;
  assign mem_MPORT_177_en = reset;
  assign mem_MPORT_178_data = 2'h0;
  assign mem_MPORT_178_addr = 8'hb2;
  assign mem_MPORT_178_mask = 1'h1;
  assign mem_MPORT_178_en = reset;
  assign mem_MPORT_179_data = 2'h0;
  assign mem_MPORT_179_addr = 8'hb3;
  assign mem_MPORT_179_mask = 1'h1;
  assign mem_MPORT_179_en = reset;
  assign mem_MPORT_180_data = 2'h0;
  assign mem_MPORT_180_addr = 8'hb4;
  assign mem_MPORT_180_mask = 1'h1;
  assign mem_MPORT_180_en = reset;
  assign mem_MPORT_181_data = 2'h0;
  assign mem_MPORT_181_addr = 8'hb5;
  assign mem_MPORT_181_mask = 1'h1;
  assign mem_MPORT_181_en = reset;
  assign mem_MPORT_182_data = 2'h0;
  assign mem_MPORT_182_addr = 8'hb6;
  assign mem_MPORT_182_mask = 1'h1;
  assign mem_MPORT_182_en = reset;
  assign mem_MPORT_183_data = 2'h0;
  assign mem_MPORT_183_addr = 8'hb7;
  assign mem_MPORT_183_mask = 1'h1;
  assign mem_MPORT_183_en = reset;
  assign mem_MPORT_184_data = 2'h0;
  assign mem_MPORT_184_addr = 8'hb8;
  assign mem_MPORT_184_mask = 1'h1;
  assign mem_MPORT_184_en = reset;
  assign mem_MPORT_185_data = 2'h0;
  assign mem_MPORT_185_addr = 8'hb9;
  assign mem_MPORT_185_mask = 1'h1;
  assign mem_MPORT_185_en = reset;
  assign mem_MPORT_186_data = 2'h0;
  assign mem_MPORT_186_addr = 8'hba;
  assign mem_MPORT_186_mask = 1'h1;
  assign mem_MPORT_186_en = reset;
  assign mem_MPORT_187_data = 2'h0;
  assign mem_MPORT_187_addr = 8'hbb;
  assign mem_MPORT_187_mask = 1'h1;
  assign mem_MPORT_187_en = reset;
  assign mem_MPORT_188_data = 2'h0;
  assign mem_MPORT_188_addr = 8'hbc;
  assign mem_MPORT_188_mask = 1'h1;
  assign mem_MPORT_188_en = reset;
  assign mem_MPORT_189_data = 2'h0;
  assign mem_MPORT_189_addr = 8'hbd;
  assign mem_MPORT_189_mask = 1'h1;
  assign mem_MPORT_189_en = reset;
  assign mem_MPORT_190_data = 2'h0;
  assign mem_MPORT_190_addr = 8'hbe;
  assign mem_MPORT_190_mask = 1'h1;
  assign mem_MPORT_190_en = reset;
  assign mem_MPORT_191_data = 2'h0;
  assign mem_MPORT_191_addr = 8'hbf;
  assign mem_MPORT_191_mask = 1'h1;
  assign mem_MPORT_191_en = reset;
  assign mem_MPORT_192_data = 2'h0;
  assign mem_MPORT_192_addr = 8'hc0;
  assign mem_MPORT_192_mask = 1'h1;
  assign mem_MPORT_192_en = reset;
  assign mem_MPORT_193_data = 2'h0;
  assign mem_MPORT_193_addr = 8'hc1;
  assign mem_MPORT_193_mask = 1'h1;
  assign mem_MPORT_193_en = reset;
  assign mem_MPORT_194_data = 2'h0;
  assign mem_MPORT_194_addr = 8'hc2;
  assign mem_MPORT_194_mask = 1'h1;
  assign mem_MPORT_194_en = reset;
  assign mem_MPORT_195_data = 2'h0;
  assign mem_MPORT_195_addr = 8'hc3;
  assign mem_MPORT_195_mask = 1'h1;
  assign mem_MPORT_195_en = reset;
  assign mem_MPORT_196_data = 2'h0;
  assign mem_MPORT_196_addr = 8'hc4;
  assign mem_MPORT_196_mask = 1'h1;
  assign mem_MPORT_196_en = reset;
  assign mem_MPORT_197_data = 2'h0;
  assign mem_MPORT_197_addr = 8'hc5;
  assign mem_MPORT_197_mask = 1'h1;
  assign mem_MPORT_197_en = reset;
  assign mem_MPORT_198_data = 2'h0;
  assign mem_MPORT_198_addr = 8'hc6;
  assign mem_MPORT_198_mask = 1'h1;
  assign mem_MPORT_198_en = reset;
  assign mem_MPORT_199_data = 2'h0;
  assign mem_MPORT_199_addr = 8'hc7;
  assign mem_MPORT_199_mask = 1'h1;
  assign mem_MPORT_199_en = reset;
  assign mem_MPORT_200_data = 2'h0;
  assign mem_MPORT_200_addr = 8'hc8;
  assign mem_MPORT_200_mask = 1'h1;
  assign mem_MPORT_200_en = reset;
  assign mem_MPORT_201_data = 2'h0;
  assign mem_MPORT_201_addr = 8'hc9;
  assign mem_MPORT_201_mask = 1'h1;
  assign mem_MPORT_201_en = reset;
  assign mem_MPORT_202_data = 2'h0;
  assign mem_MPORT_202_addr = 8'hca;
  assign mem_MPORT_202_mask = 1'h1;
  assign mem_MPORT_202_en = reset;
  assign mem_MPORT_203_data = 2'h0;
  assign mem_MPORT_203_addr = 8'hcb;
  assign mem_MPORT_203_mask = 1'h1;
  assign mem_MPORT_203_en = reset;
  assign mem_MPORT_204_data = 2'h0;
  assign mem_MPORT_204_addr = 8'hcc;
  assign mem_MPORT_204_mask = 1'h1;
  assign mem_MPORT_204_en = reset;
  assign mem_MPORT_205_data = 2'h0;
  assign mem_MPORT_205_addr = 8'hcd;
  assign mem_MPORT_205_mask = 1'h1;
  assign mem_MPORT_205_en = reset;
  assign mem_MPORT_206_data = 2'h0;
  assign mem_MPORT_206_addr = 8'hce;
  assign mem_MPORT_206_mask = 1'h1;
  assign mem_MPORT_206_en = reset;
  assign mem_MPORT_207_data = 2'h0;
  assign mem_MPORT_207_addr = 8'hcf;
  assign mem_MPORT_207_mask = 1'h1;
  assign mem_MPORT_207_en = reset;
  assign mem_MPORT_208_data = 2'h0;
  assign mem_MPORT_208_addr = 8'hd0;
  assign mem_MPORT_208_mask = 1'h1;
  assign mem_MPORT_208_en = reset;
  assign mem_MPORT_209_data = 2'h0;
  assign mem_MPORT_209_addr = 8'hd1;
  assign mem_MPORT_209_mask = 1'h1;
  assign mem_MPORT_209_en = reset;
  assign mem_MPORT_210_data = 2'h0;
  assign mem_MPORT_210_addr = 8'hd2;
  assign mem_MPORT_210_mask = 1'h1;
  assign mem_MPORT_210_en = reset;
  assign mem_MPORT_211_data = 2'h0;
  assign mem_MPORT_211_addr = 8'hd3;
  assign mem_MPORT_211_mask = 1'h1;
  assign mem_MPORT_211_en = reset;
  assign mem_MPORT_212_data = 2'h0;
  assign mem_MPORT_212_addr = 8'hd4;
  assign mem_MPORT_212_mask = 1'h1;
  assign mem_MPORT_212_en = reset;
  assign mem_MPORT_213_data = 2'h0;
  assign mem_MPORT_213_addr = 8'hd5;
  assign mem_MPORT_213_mask = 1'h1;
  assign mem_MPORT_213_en = reset;
  assign mem_MPORT_214_data = 2'h0;
  assign mem_MPORT_214_addr = 8'hd6;
  assign mem_MPORT_214_mask = 1'h1;
  assign mem_MPORT_214_en = reset;
  assign mem_MPORT_215_data = 2'h0;
  assign mem_MPORT_215_addr = 8'hd7;
  assign mem_MPORT_215_mask = 1'h1;
  assign mem_MPORT_215_en = reset;
  assign mem_MPORT_216_data = 2'h0;
  assign mem_MPORT_216_addr = 8'hd8;
  assign mem_MPORT_216_mask = 1'h1;
  assign mem_MPORT_216_en = reset;
  assign mem_MPORT_217_data = 2'h0;
  assign mem_MPORT_217_addr = 8'hd9;
  assign mem_MPORT_217_mask = 1'h1;
  assign mem_MPORT_217_en = reset;
  assign mem_MPORT_218_data = 2'h0;
  assign mem_MPORT_218_addr = 8'hda;
  assign mem_MPORT_218_mask = 1'h1;
  assign mem_MPORT_218_en = reset;
  assign mem_MPORT_219_data = 2'h0;
  assign mem_MPORT_219_addr = 8'hdb;
  assign mem_MPORT_219_mask = 1'h1;
  assign mem_MPORT_219_en = reset;
  assign mem_MPORT_220_data = 2'h0;
  assign mem_MPORT_220_addr = 8'hdc;
  assign mem_MPORT_220_mask = 1'h1;
  assign mem_MPORT_220_en = reset;
  assign mem_MPORT_221_data = 2'h0;
  assign mem_MPORT_221_addr = 8'hdd;
  assign mem_MPORT_221_mask = 1'h1;
  assign mem_MPORT_221_en = reset;
  assign mem_MPORT_222_data = 2'h0;
  assign mem_MPORT_222_addr = 8'hde;
  assign mem_MPORT_222_mask = 1'h1;
  assign mem_MPORT_222_en = reset;
  assign mem_MPORT_223_data = 2'h0;
  assign mem_MPORT_223_addr = 8'hdf;
  assign mem_MPORT_223_mask = 1'h1;
  assign mem_MPORT_223_en = reset;
  assign mem_MPORT_224_data = 2'h0;
  assign mem_MPORT_224_addr = 8'he0;
  assign mem_MPORT_224_mask = 1'h1;
  assign mem_MPORT_224_en = reset;
  assign mem_MPORT_225_data = 2'h0;
  assign mem_MPORT_225_addr = 8'he1;
  assign mem_MPORT_225_mask = 1'h1;
  assign mem_MPORT_225_en = reset;
  assign mem_MPORT_226_data = 2'h0;
  assign mem_MPORT_226_addr = 8'he2;
  assign mem_MPORT_226_mask = 1'h1;
  assign mem_MPORT_226_en = reset;
  assign mem_MPORT_227_data = 2'h0;
  assign mem_MPORT_227_addr = 8'he3;
  assign mem_MPORT_227_mask = 1'h1;
  assign mem_MPORT_227_en = reset;
  assign mem_MPORT_228_data = 2'h0;
  assign mem_MPORT_228_addr = 8'he4;
  assign mem_MPORT_228_mask = 1'h1;
  assign mem_MPORT_228_en = reset;
  assign mem_MPORT_229_data = 2'h0;
  assign mem_MPORT_229_addr = 8'he5;
  assign mem_MPORT_229_mask = 1'h1;
  assign mem_MPORT_229_en = reset;
  assign mem_MPORT_230_data = 2'h0;
  assign mem_MPORT_230_addr = 8'he6;
  assign mem_MPORT_230_mask = 1'h1;
  assign mem_MPORT_230_en = reset;
  assign mem_MPORT_231_data = 2'h0;
  assign mem_MPORT_231_addr = 8'he7;
  assign mem_MPORT_231_mask = 1'h1;
  assign mem_MPORT_231_en = reset;
  assign mem_MPORT_232_data = 2'h0;
  assign mem_MPORT_232_addr = 8'he8;
  assign mem_MPORT_232_mask = 1'h1;
  assign mem_MPORT_232_en = reset;
  assign mem_MPORT_233_data = 2'h0;
  assign mem_MPORT_233_addr = 8'he9;
  assign mem_MPORT_233_mask = 1'h1;
  assign mem_MPORT_233_en = reset;
  assign mem_MPORT_234_data = 2'h0;
  assign mem_MPORT_234_addr = 8'hea;
  assign mem_MPORT_234_mask = 1'h1;
  assign mem_MPORT_234_en = reset;
  assign mem_MPORT_235_data = 2'h0;
  assign mem_MPORT_235_addr = 8'heb;
  assign mem_MPORT_235_mask = 1'h1;
  assign mem_MPORT_235_en = reset;
  assign mem_MPORT_236_data = 2'h0;
  assign mem_MPORT_236_addr = 8'hec;
  assign mem_MPORT_236_mask = 1'h1;
  assign mem_MPORT_236_en = reset;
  assign mem_MPORT_237_data = 2'h0;
  assign mem_MPORT_237_addr = 8'hed;
  assign mem_MPORT_237_mask = 1'h1;
  assign mem_MPORT_237_en = reset;
  assign mem_MPORT_238_data = 2'h0;
  assign mem_MPORT_238_addr = 8'hee;
  assign mem_MPORT_238_mask = 1'h1;
  assign mem_MPORT_238_en = reset;
  assign mem_MPORT_239_data = 2'h0;
  assign mem_MPORT_239_addr = 8'hef;
  assign mem_MPORT_239_mask = 1'h1;
  assign mem_MPORT_239_en = reset;
  assign mem_MPORT_240_data = 2'h0;
  assign mem_MPORT_240_addr = 8'hf0;
  assign mem_MPORT_240_mask = 1'h1;
  assign mem_MPORT_240_en = reset;
  assign mem_MPORT_241_data = 2'h0;
  assign mem_MPORT_241_addr = 8'hf1;
  assign mem_MPORT_241_mask = 1'h1;
  assign mem_MPORT_241_en = reset;
  assign mem_MPORT_242_data = 2'h0;
  assign mem_MPORT_242_addr = 8'hf2;
  assign mem_MPORT_242_mask = 1'h1;
  assign mem_MPORT_242_en = reset;
  assign mem_MPORT_243_data = 2'h0;
  assign mem_MPORT_243_addr = 8'hf3;
  assign mem_MPORT_243_mask = 1'h1;
  assign mem_MPORT_243_en = reset;
  assign mem_MPORT_244_data = 2'h0;
  assign mem_MPORT_244_addr = 8'hf4;
  assign mem_MPORT_244_mask = 1'h1;
  assign mem_MPORT_244_en = reset;
  assign mem_MPORT_245_data = 2'h0;
  assign mem_MPORT_245_addr = 8'hf5;
  assign mem_MPORT_245_mask = 1'h1;
  assign mem_MPORT_245_en = reset;
  assign mem_MPORT_246_data = 2'h0;
  assign mem_MPORT_246_addr = 8'hf6;
  assign mem_MPORT_246_mask = 1'h1;
  assign mem_MPORT_246_en = reset;
  assign mem_MPORT_247_data = 2'h0;
  assign mem_MPORT_247_addr = 8'hf7;
  assign mem_MPORT_247_mask = 1'h1;
  assign mem_MPORT_247_en = reset;
  assign mem_MPORT_248_data = 2'h0;
  assign mem_MPORT_248_addr = 8'hf8;
  assign mem_MPORT_248_mask = 1'h1;
  assign mem_MPORT_248_en = reset;
  assign mem_MPORT_249_data = 2'h0;
  assign mem_MPORT_249_addr = 8'hf9;
  assign mem_MPORT_249_mask = 1'h1;
  assign mem_MPORT_249_en = reset;
  assign mem_MPORT_250_data = 2'h0;
  assign mem_MPORT_250_addr = 8'hfa;
  assign mem_MPORT_250_mask = 1'h1;
  assign mem_MPORT_250_en = reset;
  assign mem_MPORT_251_data = 2'h0;
  assign mem_MPORT_251_addr = 8'hfb;
  assign mem_MPORT_251_mask = 1'h1;
  assign mem_MPORT_251_en = reset;
  assign mem_MPORT_252_data = 2'h0;
  assign mem_MPORT_252_addr = 8'hfc;
  assign mem_MPORT_252_mask = 1'h1;
  assign mem_MPORT_252_en = reset;
  assign mem_MPORT_253_data = 2'h0;
  assign mem_MPORT_253_addr = 8'hfd;
  assign mem_MPORT_253_mask = 1'h1;
  assign mem_MPORT_253_en = reset;
  assign mem_MPORT_254_data = 2'h0;
  assign mem_MPORT_254_addr = 8'hfe;
  assign mem_MPORT_254_mask = 1'h1;
  assign mem_MPORT_254_en = reset;
  assign mem_MPORT_255_data = 2'h0;
  assign mem_MPORT_255_addr = 8'hff;
  assign mem_MPORT_255_mask = 1'h1;
  assign mem_MPORT_255_en = reset;
  assign mem_MPORT_256_data = io_w_data;
  assign mem_MPORT_256_addr = io_w_addr;
  assign mem_MPORT_256_mask = 1'h1;
  assign mem_MPORT_256_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_129_en & mem_MPORT_129_mask) begin
      mem[mem_MPORT_129_addr] <= mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_130_en & mem_MPORT_130_mask) begin
      mem[mem_MPORT_130_addr] <= mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_131_en & mem_MPORT_131_mask) begin
      mem[mem_MPORT_131_addr] <= mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_132_en & mem_MPORT_132_mask) begin
      mem[mem_MPORT_132_addr] <= mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_133_en & mem_MPORT_133_mask) begin
      mem[mem_MPORT_133_addr] <= mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_134_en & mem_MPORT_134_mask) begin
      mem[mem_MPORT_134_addr] <= mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_135_en & mem_MPORT_135_mask) begin
      mem[mem_MPORT_135_addr] <= mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_136_en & mem_MPORT_136_mask) begin
      mem[mem_MPORT_136_addr] <= mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_137_en & mem_MPORT_137_mask) begin
      mem[mem_MPORT_137_addr] <= mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_138_en & mem_MPORT_138_mask) begin
      mem[mem_MPORT_138_addr] <= mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_139_en & mem_MPORT_139_mask) begin
      mem[mem_MPORT_139_addr] <= mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_140_en & mem_MPORT_140_mask) begin
      mem[mem_MPORT_140_addr] <= mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_141_en & mem_MPORT_141_mask) begin
      mem[mem_MPORT_141_addr] <= mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_142_en & mem_MPORT_142_mask) begin
      mem[mem_MPORT_142_addr] <= mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_143_en & mem_MPORT_143_mask) begin
      mem[mem_MPORT_143_addr] <= mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_144_en & mem_MPORT_144_mask) begin
      mem[mem_MPORT_144_addr] <= mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_145_en & mem_MPORT_145_mask) begin
      mem[mem_MPORT_145_addr] <= mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_146_en & mem_MPORT_146_mask) begin
      mem[mem_MPORT_146_addr] <= mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_147_en & mem_MPORT_147_mask) begin
      mem[mem_MPORT_147_addr] <= mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_148_en & mem_MPORT_148_mask) begin
      mem[mem_MPORT_148_addr] <= mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_149_en & mem_MPORT_149_mask) begin
      mem[mem_MPORT_149_addr] <= mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_150_en & mem_MPORT_150_mask) begin
      mem[mem_MPORT_150_addr] <= mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_151_en & mem_MPORT_151_mask) begin
      mem[mem_MPORT_151_addr] <= mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_152_en & mem_MPORT_152_mask) begin
      mem[mem_MPORT_152_addr] <= mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_153_en & mem_MPORT_153_mask) begin
      mem[mem_MPORT_153_addr] <= mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_154_en & mem_MPORT_154_mask) begin
      mem[mem_MPORT_154_addr] <= mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_155_en & mem_MPORT_155_mask) begin
      mem[mem_MPORT_155_addr] <= mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_156_en & mem_MPORT_156_mask) begin
      mem[mem_MPORT_156_addr] <= mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_157_en & mem_MPORT_157_mask) begin
      mem[mem_MPORT_157_addr] <= mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_158_en & mem_MPORT_158_mask) begin
      mem[mem_MPORT_158_addr] <= mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_159_en & mem_MPORT_159_mask) begin
      mem[mem_MPORT_159_addr] <= mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_160_en & mem_MPORT_160_mask) begin
      mem[mem_MPORT_160_addr] <= mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_161_en & mem_MPORT_161_mask) begin
      mem[mem_MPORT_161_addr] <= mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_162_en & mem_MPORT_162_mask) begin
      mem[mem_MPORT_162_addr] <= mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_163_en & mem_MPORT_163_mask) begin
      mem[mem_MPORT_163_addr] <= mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_164_en & mem_MPORT_164_mask) begin
      mem[mem_MPORT_164_addr] <= mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_165_en & mem_MPORT_165_mask) begin
      mem[mem_MPORT_165_addr] <= mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_166_en & mem_MPORT_166_mask) begin
      mem[mem_MPORT_166_addr] <= mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_167_en & mem_MPORT_167_mask) begin
      mem[mem_MPORT_167_addr] <= mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_168_en & mem_MPORT_168_mask) begin
      mem[mem_MPORT_168_addr] <= mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_169_en & mem_MPORT_169_mask) begin
      mem[mem_MPORT_169_addr] <= mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_170_en & mem_MPORT_170_mask) begin
      mem[mem_MPORT_170_addr] <= mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_171_en & mem_MPORT_171_mask) begin
      mem[mem_MPORT_171_addr] <= mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_172_en & mem_MPORT_172_mask) begin
      mem[mem_MPORT_172_addr] <= mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_173_en & mem_MPORT_173_mask) begin
      mem[mem_MPORT_173_addr] <= mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_174_en & mem_MPORT_174_mask) begin
      mem[mem_MPORT_174_addr] <= mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_175_en & mem_MPORT_175_mask) begin
      mem[mem_MPORT_175_addr] <= mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_176_en & mem_MPORT_176_mask) begin
      mem[mem_MPORT_176_addr] <= mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_177_en & mem_MPORT_177_mask) begin
      mem[mem_MPORT_177_addr] <= mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_178_en & mem_MPORT_178_mask) begin
      mem[mem_MPORT_178_addr] <= mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_179_en & mem_MPORT_179_mask) begin
      mem[mem_MPORT_179_addr] <= mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_180_en & mem_MPORT_180_mask) begin
      mem[mem_MPORT_180_addr] <= mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_181_en & mem_MPORT_181_mask) begin
      mem[mem_MPORT_181_addr] <= mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_182_en & mem_MPORT_182_mask) begin
      mem[mem_MPORT_182_addr] <= mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_183_en & mem_MPORT_183_mask) begin
      mem[mem_MPORT_183_addr] <= mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_184_en & mem_MPORT_184_mask) begin
      mem[mem_MPORT_184_addr] <= mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_185_en & mem_MPORT_185_mask) begin
      mem[mem_MPORT_185_addr] <= mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_186_en & mem_MPORT_186_mask) begin
      mem[mem_MPORT_186_addr] <= mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_187_en & mem_MPORT_187_mask) begin
      mem[mem_MPORT_187_addr] <= mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_188_en & mem_MPORT_188_mask) begin
      mem[mem_MPORT_188_addr] <= mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_189_en & mem_MPORT_189_mask) begin
      mem[mem_MPORT_189_addr] <= mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_190_en & mem_MPORT_190_mask) begin
      mem[mem_MPORT_190_addr] <= mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_191_en & mem_MPORT_191_mask) begin
      mem[mem_MPORT_191_addr] <= mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_192_en & mem_MPORT_192_mask) begin
      mem[mem_MPORT_192_addr] <= mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_193_en & mem_MPORT_193_mask) begin
      mem[mem_MPORT_193_addr] <= mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_194_en & mem_MPORT_194_mask) begin
      mem[mem_MPORT_194_addr] <= mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_195_en & mem_MPORT_195_mask) begin
      mem[mem_MPORT_195_addr] <= mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_196_en & mem_MPORT_196_mask) begin
      mem[mem_MPORT_196_addr] <= mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_197_en & mem_MPORT_197_mask) begin
      mem[mem_MPORT_197_addr] <= mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_198_en & mem_MPORT_198_mask) begin
      mem[mem_MPORT_198_addr] <= mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_199_en & mem_MPORT_199_mask) begin
      mem[mem_MPORT_199_addr] <= mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_200_en & mem_MPORT_200_mask) begin
      mem[mem_MPORT_200_addr] <= mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_201_en & mem_MPORT_201_mask) begin
      mem[mem_MPORT_201_addr] <= mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_202_en & mem_MPORT_202_mask) begin
      mem[mem_MPORT_202_addr] <= mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_203_en & mem_MPORT_203_mask) begin
      mem[mem_MPORT_203_addr] <= mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_204_en & mem_MPORT_204_mask) begin
      mem[mem_MPORT_204_addr] <= mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_205_en & mem_MPORT_205_mask) begin
      mem[mem_MPORT_205_addr] <= mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_206_en & mem_MPORT_206_mask) begin
      mem[mem_MPORT_206_addr] <= mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_207_en & mem_MPORT_207_mask) begin
      mem[mem_MPORT_207_addr] <= mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_208_en & mem_MPORT_208_mask) begin
      mem[mem_MPORT_208_addr] <= mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_209_en & mem_MPORT_209_mask) begin
      mem[mem_MPORT_209_addr] <= mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_210_en & mem_MPORT_210_mask) begin
      mem[mem_MPORT_210_addr] <= mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_211_en & mem_MPORT_211_mask) begin
      mem[mem_MPORT_211_addr] <= mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_212_en & mem_MPORT_212_mask) begin
      mem[mem_MPORT_212_addr] <= mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_213_en & mem_MPORT_213_mask) begin
      mem[mem_MPORT_213_addr] <= mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_214_en & mem_MPORT_214_mask) begin
      mem[mem_MPORT_214_addr] <= mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_215_en & mem_MPORT_215_mask) begin
      mem[mem_MPORT_215_addr] <= mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_216_en & mem_MPORT_216_mask) begin
      mem[mem_MPORT_216_addr] <= mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_217_en & mem_MPORT_217_mask) begin
      mem[mem_MPORT_217_addr] <= mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_218_en & mem_MPORT_218_mask) begin
      mem[mem_MPORT_218_addr] <= mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_219_en & mem_MPORT_219_mask) begin
      mem[mem_MPORT_219_addr] <= mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_220_en & mem_MPORT_220_mask) begin
      mem[mem_MPORT_220_addr] <= mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_221_en & mem_MPORT_221_mask) begin
      mem[mem_MPORT_221_addr] <= mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_222_en & mem_MPORT_222_mask) begin
      mem[mem_MPORT_222_addr] <= mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_223_en & mem_MPORT_223_mask) begin
      mem[mem_MPORT_223_addr] <= mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_224_en & mem_MPORT_224_mask) begin
      mem[mem_MPORT_224_addr] <= mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_225_en & mem_MPORT_225_mask) begin
      mem[mem_MPORT_225_addr] <= mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_226_en & mem_MPORT_226_mask) begin
      mem[mem_MPORT_226_addr] <= mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_227_en & mem_MPORT_227_mask) begin
      mem[mem_MPORT_227_addr] <= mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_228_en & mem_MPORT_228_mask) begin
      mem[mem_MPORT_228_addr] <= mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_229_en & mem_MPORT_229_mask) begin
      mem[mem_MPORT_229_addr] <= mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_230_en & mem_MPORT_230_mask) begin
      mem[mem_MPORT_230_addr] <= mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_231_en & mem_MPORT_231_mask) begin
      mem[mem_MPORT_231_addr] <= mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_232_en & mem_MPORT_232_mask) begin
      mem[mem_MPORT_232_addr] <= mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_233_en & mem_MPORT_233_mask) begin
      mem[mem_MPORT_233_addr] <= mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_234_en & mem_MPORT_234_mask) begin
      mem[mem_MPORT_234_addr] <= mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_235_en & mem_MPORT_235_mask) begin
      mem[mem_MPORT_235_addr] <= mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_236_en & mem_MPORT_236_mask) begin
      mem[mem_MPORT_236_addr] <= mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_237_en & mem_MPORT_237_mask) begin
      mem[mem_MPORT_237_addr] <= mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_238_en & mem_MPORT_238_mask) begin
      mem[mem_MPORT_238_addr] <= mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_239_en & mem_MPORT_239_mask) begin
      mem[mem_MPORT_239_addr] <= mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_240_en & mem_MPORT_240_mask) begin
      mem[mem_MPORT_240_addr] <= mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_241_en & mem_MPORT_241_mask) begin
      mem[mem_MPORT_241_addr] <= mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_242_en & mem_MPORT_242_mask) begin
      mem[mem_MPORT_242_addr] <= mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_243_en & mem_MPORT_243_mask) begin
      mem[mem_MPORT_243_addr] <= mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_244_en & mem_MPORT_244_mask) begin
      mem[mem_MPORT_244_addr] <= mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_245_en & mem_MPORT_245_mask) begin
      mem[mem_MPORT_245_addr] <= mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_246_en & mem_MPORT_246_mask) begin
      mem[mem_MPORT_246_addr] <= mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_247_en & mem_MPORT_247_mask) begin
      mem[mem_MPORT_247_addr] <= mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_248_en & mem_MPORT_248_mask) begin
      mem[mem_MPORT_248_addr] <= mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_249_en & mem_MPORT_249_mask) begin
      mem[mem_MPORT_249_addr] <= mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_250_en & mem_MPORT_250_mask) begin
      mem[mem_MPORT_250_addr] <= mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_251_en & mem_MPORT_251_mask) begin
      mem[mem_MPORT_251_addr] <= mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_252_en & mem_MPORT_252_mask) begin
      mem[mem_MPORT_252_addr] <= mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_253_en & mem_MPORT_253_mask) begin
      mem[mem_MPORT_253_addr] <= mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_254_en & mem_MPORT_254_mask) begin
      mem[mem_MPORT_254_addr] <= mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_255_en & mem_MPORT_255_mask) begin
      mem[mem_MPORT_255_addr] <= mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_256_en & mem_MPORT_256_mask) begin
      mem[mem_MPORT_256_addr] <= mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMArray_2P_19(
  input        clock,
  input        reset,
  input  [7:0] io_r_addr,
  output [1:0] io_r_data_0,
  output [1:0] io_r_data_1,
  output [1:0] io_r_data_2,
  output [1:0] io_r_data_3,
  output [1:0] io_r_data_4,
  output [1:0] io_r_data_5,
  output [1:0] io_r_data_6,
  output [1:0] io_r_data_7,
  input        io_w_en,
  input  [7:0] io_w_addr,
  input  [1:0] io_w_data_0,
  input  [1:0] io_w_data_1,
  input  [1:0] io_w_data_2,
  input  [1:0] io_w_data_3,
  input  [1:0] io_w_data_4,
  input  [1:0] io_w_data_5,
  input  [1:0] io_w_data_6,
  input  [1:0] io_w_data_7,
  input  [7:0] io_w_maskOH
);
  wire  brams_0_clock; // @[SRAM_1.scala 201:38]
  wire  brams_0_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_0_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_0_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_0_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_0_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_0_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_clock; // @[SRAM_1.scala 201:38]
  wire  brams_1_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_1_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_1_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_1_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_1_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_1_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_clock; // @[SRAM_1.scala 201:38]
  wire  brams_2_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_2_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_2_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_2_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_2_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_2_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_clock; // @[SRAM_1.scala 201:38]
  wire  brams_3_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_3_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_3_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_3_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_3_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_3_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_clock; // @[SRAM_1.scala 201:38]
  wire  brams_4_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_4_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_4_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_4_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_4_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_4_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_clock; // @[SRAM_1.scala 201:38]
  wire  brams_5_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_5_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_5_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_5_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_5_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_5_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_clock; // @[SRAM_1.scala 201:38]
  wire  brams_6_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_6_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_6_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_6_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_6_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_6_io_w_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_clock; // @[SRAM_1.scala 201:38]
  wire  brams_7_reset; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_7_io_r_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_7_io_r_data; // @[SRAM_1.scala 201:38]
  wire  brams_7_io_w_en; // @[SRAM_1.scala 201:38]
  wire [7:0] brams_7_io_w_addr; // @[SRAM_1.scala 201:38]
  wire [1:0] brams_7_io_w_data; // @[SRAM_1.scala 201:38]
  BankRAM_2P_120 brams_0 ( // @[SRAM_1.scala 201:38]
    .clock(brams_0_clock),
    .reset(brams_0_reset),
    .io_r_addr(brams_0_io_r_addr),
    .io_r_data(brams_0_io_r_data),
    .io_w_en(brams_0_io_w_en),
    .io_w_addr(brams_0_io_w_addr),
    .io_w_data(brams_0_io_w_data)
  );
  BankRAM_2P_120 brams_1 ( // @[SRAM_1.scala 201:38]
    .clock(brams_1_clock),
    .reset(brams_1_reset),
    .io_r_addr(brams_1_io_r_addr),
    .io_r_data(brams_1_io_r_data),
    .io_w_en(brams_1_io_w_en),
    .io_w_addr(brams_1_io_w_addr),
    .io_w_data(brams_1_io_w_data)
  );
  BankRAM_2P_120 brams_2 ( // @[SRAM_1.scala 201:38]
    .clock(brams_2_clock),
    .reset(brams_2_reset),
    .io_r_addr(brams_2_io_r_addr),
    .io_r_data(brams_2_io_r_data),
    .io_w_en(brams_2_io_w_en),
    .io_w_addr(brams_2_io_w_addr),
    .io_w_data(brams_2_io_w_data)
  );
  BankRAM_2P_120 brams_3 ( // @[SRAM_1.scala 201:38]
    .clock(brams_3_clock),
    .reset(brams_3_reset),
    .io_r_addr(brams_3_io_r_addr),
    .io_r_data(brams_3_io_r_data),
    .io_w_en(brams_3_io_w_en),
    .io_w_addr(brams_3_io_w_addr),
    .io_w_data(brams_3_io_w_data)
  );
  BankRAM_2P_120 brams_4 ( // @[SRAM_1.scala 201:38]
    .clock(brams_4_clock),
    .reset(brams_4_reset),
    .io_r_addr(brams_4_io_r_addr),
    .io_r_data(brams_4_io_r_data),
    .io_w_en(brams_4_io_w_en),
    .io_w_addr(brams_4_io_w_addr),
    .io_w_data(brams_4_io_w_data)
  );
  BankRAM_2P_120 brams_5 ( // @[SRAM_1.scala 201:38]
    .clock(brams_5_clock),
    .reset(brams_5_reset),
    .io_r_addr(brams_5_io_r_addr),
    .io_r_data(brams_5_io_r_data),
    .io_w_en(brams_5_io_w_en),
    .io_w_addr(brams_5_io_w_addr),
    .io_w_data(brams_5_io_w_data)
  );
  BankRAM_2P_120 brams_6 ( // @[SRAM_1.scala 201:38]
    .clock(brams_6_clock),
    .reset(brams_6_reset),
    .io_r_addr(brams_6_io_r_addr),
    .io_r_data(brams_6_io_r_data),
    .io_w_en(brams_6_io_w_en),
    .io_w_addr(brams_6_io_w_addr),
    .io_w_data(brams_6_io_w_data)
  );
  BankRAM_2P_120 brams_7 ( // @[SRAM_1.scala 201:38]
    .clock(brams_7_clock),
    .reset(brams_7_reset),
    .io_r_addr(brams_7_io_r_addr),
    .io_r_data(brams_7_io_r_data),
    .io_w_en(brams_7_io_w_en),
    .io_w_addr(brams_7_io_w_addr),
    .io_w_data(brams_7_io_w_data)
  );
  assign io_r_data_0 = brams_0_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_1 = brams_1_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_2 = brams_2_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_3 = brams_3_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_4 = brams_4_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_5 = brams_5_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_6 = brams_6_io_r_data; // @[SRAM_1.scala 206:22]
  assign io_r_data_7 = brams_7_io_r_data; // @[SRAM_1.scala 206:22]
  assign brams_0_clock = clock;
  assign brams_0_reset = reset;
  assign brams_0_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_0_io_w_en = io_w_en & io_w_maskOH[0]; // @[SRAM_1.scala 208:37]
  assign brams_0_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_0_io_w_data = io_w_data_0; // @[SRAM_1.scala 210:28]
  assign brams_1_clock = clock;
  assign brams_1_reset = reset;
  assign brams_1_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_1_io_w_en = io_w_en & io_w_maskOH[1]; // @[SRAM_1.scala 208:37]
  assign brams_1_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_1_io_w_data = io_w_data_1; // @[SRAM_1.scala 210:28]
  assign brams_2_clock = clock;
  assign brams_2_reset = reset;
  assign brams_2_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_2_io_w_en = io_w_en & io_w_maskOH[2]; // @[SRAM_1.scala 208:37]
  assign brams_2_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_2_io_w_data = io_w_data_2; // @[SRAM_1.scala 210:28]
  assign brams_3_clock = clock;
  assign brams_3_reset = reset;
  assign brams_3_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_3_io_w_en = io_w_en & io_w_maskOH[3]; // @[SRAM_1.scala 208:37]
  assign brams_3_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_3_io_w_data = io_w_data_3; // @[SRAM_1.scala 210:28]
  assign brams_4_clock = clock;
  assign brams_4_reset = reset;
  assign brams_4_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_4_io_w_en = io_w_en & io_w_maskOH[4]; // @[SRAM_1.scala 208:37]
  assign brams_4_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_4_io_w_data = io_w_data_4; // @[SRAM_1.scala 210:28]
  assign brams_5_clock = clock;
  assign brams_5_reset = reset;
  assign brams_5_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_5_io_w_en = io_w_en & io_w_maskOH[5]; // @[SRAM_1.scala 208:37]
  assign brams_5_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_5_io_w_data = io_w_data_5; // @[SRAM_1.scala 210:28]
  assign brams_6_clock = clock;
  assign brams_6_reset = reset;
  assign brams_6_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_6_io_w_en = io_w_en & io_w_maskOH[6]; // @[SRAM_1.scala 208:37]
  assign brams_6_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_6_io_w_data = io_w_data_6; // @[SRAM_1.scala 210:28]
  assign brams_7_clock = clock;
  assign brams_7_reset = reset;
  assign brams_7_io_r_addr = io_r_addr; // @[SRAM_1.scala 205:28]
  assign brams_7_io_w_en = io_w_en & io_w_maskOH[7]; // @[SRAM_1.scala 208:37]
  assign brams_7_io_w_addr = io_w_addr; // @[SRAM_1.scala 209:28]
  assign brams_7_io_w_data = io_w_data_7; // @[SRAM_1.scala 210:28]
endmodule
module DCacheDirectory_1(
  input         clock,
  input         reset,
  output        io_read_req_ready,
  input         io_read_req_valid,
  input  [31:0] io_read_req_bits_addr,
  output        io_read_resp_bits_hit,
  output [7:0]  io_read_resp_bits_chosenWay,
  output        io_read_resp_bits_isDirtyWay,
  output [19:0] io_read_resp_bits_tagRdVec_0,
  output [19:0] io_read_resp_bits_tagRdVec_1,
  output [19:0] io_read_resp_bits_tagRdVec_2,
  output [19:0] io_read_resp_bits_tagRdVec_3,
  output [19:0] io_read_resp_bits_tagRdVec_4,
  output [19:0] io_read_resp_bits_tagRdVec_5,
  output [19:0] io_read_resp_bits_tagRdVec_6,
  output [19:0] io_read_resp_bits_tagRdVec_7,
  output        io_write_req_ready,
  input         io_write_req_valid,
  input  [31:0] io_write_req_bits_addr,
  input  [7:0]  io_write_req_bits_way,
  input  [1:0]  io_write_req_bits_meta
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  tagArray_clock; // @[SRAM_1.scala 255:31]
  wire  tagArray_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] tagArray_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  tagArray_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] tagArray_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [19:0] tagArray_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] tagArray_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  metaArray_clock; // @[SRAM_1.scala 255:31]
  wire  metaArray_reset; // @[SRAM_1.scala 255:31]
  wire [7:0] metaArray_io_r_addr; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_0; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_1; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_2; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_3; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_4; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_5; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_6; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_r_data_7; // @[SRAM_1.scala 255:31]
  wire  metaArray_io_w_en; // @[SRAM_1.scala 255:31]
  wire [7:0] metaArray_io_w_addr; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_0; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_1; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_2; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_3; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_4; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_5; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_6; // @[SRAM_1.scala 255:31]
  wire [1:0] metaArray_io_w_data_7; // @[SRAM_1.scala 255:31]
  wire [7:0] metaArray_io_w_maskOH; // @[SRAM_1.scala 255:31]
  wire  replaceWay_lfsr_prng_clock; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_reset; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  replaceWay_lfsr_prng_io_out_15; // @[PRNG.scala 91:22]
  wire [7:0] rSet = io_read_req_bits_addr[11:4]; // @[Parameters.scala 50:11]
  wire [19:0] rTag = io_read_req_bits_addr[31:12]; // @[Parameters.scala 46:11]
  wire  ren = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  wire [7:0] wSet = io_write_req_bits_addr[11:4]; // @[Parameters.scala 50:11]
  wire [19:0] wTag = io_write_req_bits_addr[31:12]; // @[Parameters.scala 46:11]
  wire  wen = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _T_8 = io_write_req_bits_way[0] + io_write_req_bits_way[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_10 = io_write_req_bits_way[2] + io_write_req_bits_way[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_12 = _T_8 + _T_10; // @[Bitwise.scala 51:90]
  wire [1:0] _T_14 = io_write_req_bits_way[4] + io_write_req_bits_way[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_16 = io_write_req_bits_way[6] + io_write_req_bits_way[7]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_18 = _T_14 + _T_16; // @[Bitwise.scala 51:90]
  wire [3:0] _T_20 = _T_12 + _T_18; // @[Bitwise.scala 51:90]
  wire  _T_46 = ~reset; // @[Directory.scala 69:11]
  wire [19:0] rdata__0 = ren ? tagArray_io_r_data_0 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__1 = ren ? tagArray_io_r_data_1 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__2 = ren ? tagArray_io_r_data_2 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__3 = ren ? tagArray_io_r_data_3 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__4 = ren ? tagArray_io_r_data_4 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__5 = ren ? tagArray_io_r_data_5 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__6 = ren ? tagArray_io_r_data_6 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [19:0] rdata__7 = ren ? tagArray_io_r_data_7 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_0 = ren ? metaArray_io_r_data_0 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_1 = ren ? metaArray_io_r_data_1 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_2 = ren ? metaArray_io_r_data_2 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_3 = ren ? metaArray_io_r_data_3 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_4 = ren ? metaArray_io_r_data_4 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_5 = ren ? metaArray_io_r_data_5 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_6 = ren ? metaArray_io_r_data_6 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [1:0] rdata_1_7 = ren ? metaArray_io_r_data_7 : 2'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  wire [15:0] _T_48 = {rdata_1_7,rdata_1_6,rdata_1_5,rdata_1_4,rdata_1_3,rdata_1_2,rdata_1_1,rdata_1_0}; // @[Directory.scala 82:52]
  wire  metaRdVec_0_valid = _T_48[0]; // @[Directory.scala 82:52]
  wire  metaRdVec_0_dirty = _T_48[1]; // @[Directory.scala 82:52]
  wire  metaRdVec_1_valid = _T_48[2]; // @[Directory.scala 82:52]
  wire  metaRdVec_1_dirty = _T_48[3]; // @[Directory.scala 82:52]
  wire  metaRdVec_2_valid = _T_48[4]; // @[Directory.scala 82:52]
  wire  metaRdVec_2_dirty = _T_48[5]; // @[Directory.scala 82:52]
  wire  metaRdVec_3_valid = _T_48[6]; // @[Directory.scala 82:52]
  wire  metaRdVec_3_dirty = _T_48[7]; // @[Directory.scala 82:52]
  wire  metaRdVec_4_valid = _T_48[8]; // @[Directory.scala 82:52]
  wire  metaRdVec_4_dirty = _T_48[9]; // @[Directory.scala 82:52]
  wire  metaRdVec_5_valid = _T_48[10]; // @[Directory.scala 82:52]
  wire  metaRdVec_5_dirty = _T_48[11]; // @[Directory.scala 82:52]
  wire  metaRdVec_6_valid = _T_48[12]; // @[Directory.scala 82:52]
  wire  metaRdVec_6_dirty = _T_48[13]; // @[Directory.scala 82:52]
  wire  metaRdVec_7_valid = _T_48[14]; // @[Directory.scala 82:52]
  wire  metaRdVec_7_dirty = _T_48[15]; // @[Directory.scala 82:52]
  wire  tagMatchVec_0 = rdata__0 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_1 = rdata__1 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_2 = rdata__2 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_3 = rdata__3 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_4 = rdata__4 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_5 = rdata__5 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_6 = rdata__6 == rTag; // @[Directory.scala 85:46]
  wire  tagMatchVec_7 = rdata__7 == rTag; // @[Directory.scala 85:46]
  wire  _matchWayOH_T = tagMatchVec_0 & metaRdVec_0_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_1 = tagMatchVec_1 & metaRdVec_1_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_2 = tagMatchVec_2 & metaRdVec_2_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_3 = tagMatchVec_3 & metaRdVec_3_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_4 = tagMatchVec_4 & metaRdVec_4_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_5 = tagMatchVec_5 & metaRdVec_5_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_6 = tagMatchVec_6 & metaRdVec_6_valid; // @[Directory.scala 88:80]
  wire  _matchWayOH_T_7 = tagMatchVec_7 & metaRdVec_7_valid; // @[Directory.scala 88:80]
  wire [7:0] matchWayOH = {_matchWayOH_T_7,_matchWayOH_T_6,_matchWayOH_T_5,_matchWayOH_T_4,_matchWayOH_T_3,
    _matchWayOH_T_2,_matchWayOH_T_1,_matchWayOH_T}; // @[Cat.scala 33:92]
  wire  invalidWayVec_0 = ~metaRdVec_0_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_1 = ~metaRdVec_1_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_2 = ~metaRdVec_2_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_3 = ~metaRdVec_3_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_4 = ~metaRdVec_4_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_5 = ~metaRdVec_5_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_6 = ~metaRdVec_6_valid; // @[Directory.scala 89:53]
  wire  invalidWayVec_7 = ~metaRdVec_7_valid; // @[Directory.scala 89:53]
  wire [7:0] _invalidWayOH_T_16 = invalidWayVec_6 ? 8'h40 : 8'h80; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_17 = invalidWayVec_5 ? 8'h20 : _invalidWayOH_T_16; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_18 = invalidWayVec_4 ? 8'h10 : _invalidWayOH_T_17; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_19 = invalidWayVec_3 ? 8'h8 : _invalidWayOH_T_18; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_20 = invalidWayVec_2 ? 8'h4 : _invalidWayOH_T_19; // @[Mux.scala 47:70]
  wire [7:0] _invalidWayOH_T_21 = invalidWayVec_1 ? 8'h2 : _invalidWayOH_T_20; // @[Mux.scala 47:70]
  wire [7:0] invalidWayOH = invalidWayVec_0 ? 8'h1 : _invalidWayOH_T_21; // @[Mux.scala 47:70]
  wire [7:0] _hasInvalidWay_T = {invalidWayVec_0,invalidWayVec_1,invalidWayVec_2,invalidWayVec_3,invalidWayVec_4,
    invalidWayVec_5,invalidWayVec_6,invalidWayVec_7}; // @[Cat.scala 33:92]
  wire  hasInvalidWay = |_hasInvalidWay_T; // @[Directory.scala 91:44]
  wire [7:0] replaceWay_lfsr_lo = {replaceWay_lfsr_prng_io_out_7,replaceWay_lfsr_prng_io_out_6,
    replaceWay_lfsr_prng_io_out_5,replaceWay_lfsr_prng_io_out_4,replaceWay_lfsr_prng_io_out_3,
    replaceWay_lfsr_prng_io_out_2,replaceWay_lfsr_prng_io_out_1,replaceWay_lfsr_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [15:0] replaceWay_lfsr = {replaceWay_lfsr_prng_io_out_15,replaceWay_lfsr_prng_io_out_14,
    replaceWay_lfsr_prng_io_out_13,replaceWay_lfsr_prng_io_out_12,replaceWay_lfsr_prng_io_out_11,
    replaceWay_lfsr_prng_io_out_10,replaceWay_lfsr_prng_io_out_9,replaceWay_lfsr_prng_io_out_8,replaceWay_lfsr_lo}; // @[PRNG.scala 95:17]
  wire [2:0] replaceWay_outputWay_shiftAmount = replaceWay_lfsr[2:0]; // @[DCache.scala 60:39]
  wire [7:0] replaceWay = 8'h1 << replaceWay_outputWay_shiftAmount; // @[OneHot.scala 64:12]
  wire  _replaceWayReg_T = ~io_read_req_valid; // @[Directory.scala 93:65]
  reg [7:0] replaceWayReg; // @[Reg.scala 19:16]
  wire  isHit = |matchWayOH; // @[Directory.scala 95:41]
  wire [7:0] _choseWayOH_T = hasInvalidWay ? invalidWayOH : replaceWayReg; // @[Directory.scala 96:51]
  wire [7:0] choseWayOH = isHit ? matchWayOH : _choseWayOH_T; // @[Directory.scala 96:28]
  wire [7:0] dirtyWayOH = {metaRdVec_7_dirty,metaRdVec_6_dirty,metaRdVec_5_dirty,metaRdVec_4_dirty,metaRdVec_3_dirty,
    metaRdVec_2_dirty,metaRdVec_1_dirty,metaRdVec_0_dirty}; // @[Cat.scala 33:92]
  wire [7:0] _isDirtyWay_T = choseWayOH & dirtyWayOH; // @[Directory.scala 98:38]
  wire [1:0] _T_73 = choseWayOH[0] + choseWayOH[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_75 = choseWayOH[2] + choseWayOH[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_77 = _T_73 + _T_75; // @[Bitwise.scala 51:90]
  wire [1:0] _T_79 = choseWayOH[4] + choseWayOH[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_81 = choseWayOH[6] + choseWayOH[7]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_83 = _T_79 + _T_81; // @[Bitwise.scala 51:90]
  wire [3:0] _T_85 = _T_77 + _T_83; // @[Bitwise.scala 51:90]
  SRAMArray_2P_18 tagArray ( // @[SRAM_1.scala 255:31]
    .clock(tagArray_clock),
    .reset(tagArray_reset),
    .io_r_addr(tagArray_io_r_addr),
    .io_r_data_0(tagArray_io_r_data_0),
    .io_r_data_1(tagArray_io_r_data_1),
    .io_r_data_2(tagArray_io_r_data_2),
    .io_r_data_3(tagArray_io_r_data_3),
    .io_r_data_4(tagArray_io_r_data_4),
    .io_r_data_5(tagArray_io_r_data_5),
    .io_r_data_6(tagArray_io_r_data_6),
    .io_r_data_7(tagArray_io_r_data_7),
    .io_w_en(tagArray_io_w_en),
    .io_w_addr(tagArray_io_w_addr),
    .io_w_data_0(tagArray_io_w_data_0),
    .io_w_data_1(tagArray_io_w_data_1),
    .io_w_data_2(tagArray_io_w_data_2),
    .io_w_data_3(tagArray_io_w_data_3),
    .io_w_data_4(tagArray_io_w_data_4),
    .io_w_data_5(tagArray_io_w_data_5),
    .io_w_data_6(tagArray_io_w_data_6),
    .io_w_data_7(tagArray_io_w_data_7),
    .io_w_maskOH(tagArray_io_w_maskOH)
  );
  SRAMArray_2P_19 metaArray ( // @[SRAM_1.scala 255:31]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_addr(metaArray_io_r_addr),
    .io_r_data_0(metaArray_io_r_data_0),
    .io_r_data_1(metaArray_io_r_data_1),
    .io_r_data_2(metaArray_io_r_data_2),
    .io_r_data_3(metaArray_io_r_data_3),
    .io_r_data_4(metaArray_io_r_data_4),
    .io_r_data_5(metaArray_io_r_data_5),
    .io_r_data_6(metaArray_io_r_data_6),
    .io_r_data_7(metaArray_io_r_data_7),
    .io_w_en(metaArray_io_w_en),
    .io_w_addr(metaArray_io_w_addr),
    .io_w_data_0(metaArray_io_w_data_0),
    .io_w_data_1(metaArray_io_w_data_1),
    .io_w_data_2(metaArray_io_w_data_2),
    .io_w_data_3(metaArray_io_w_data_3),
    .io_w_data_4(metaArray_io_w_data_4),
    .io_w_data_5(metaArray_io_w_data_5),
    .io_w_data_6(metaArray_io_w_data_6),
    .io_w_data_7(metaArray_io_w_data_7),
    .io_w_maskOH(metaArray_io_w_maskOH)
  );
  MaxPeriodFibonacciLFSR replaceWay_lfsr_prng ( // @[PRNG.scala 91:22]
    .clock(replaceWay_lfsr_prng_clock),
    .reset(replaceWay_lfsr_prng_reset),
    .io_out_0(replaceWay_lfsr_prng_io_out_0),
    .io_out_1(replaceWay_lfsr_prng_io_out_1),
    .io_out_2(replaceWay_lfsr_prng_io_out_2),
    .io_out_3(replaceWay_lfsr_prng_io_out_3),
    .io_out_4(replaceWay_lfsr_prng_io_out_4),
    .io_out_5(replaceWay_lfsr_prng_io_out_5),
    .io_out_6(replaceWay_lfsr_prng_io_out_6),
    .io_out_7(replaceWay_lfsr_prng_io_out_7),
    .io_out_8(replaceWay_lfsr_prng_io_out_8),
    .io_out_9(replaceWay_lfsr_prng_io_out_9),
    .io_out_10(replaceWay_lfsr_prng_io_out_10),
    .io_out_11(replaceWay_lfsr_prng_io_out_11),
    .io_out_12(replaceWay_lfsr_prng_io_out_12),
    .io_out_13(replaceWay_lfsr_prng_io_out_13),
    .io_out_14(replaceWay_lfsr_prng_io_out_14),
    .io_out_15(replaceWay_lfsr_prng_io_out_15)
  );
  assign io_read_req_ready = 1'h1; // @[Directory.scala 75:29]
  assign io_read_resp_bits_hit = |matchWayOH; // @[Directory.scala 95:41]
  assign io_read_resp_bits_chosenWay = isHit ? matchWayOH : _choseWayOH_T; // @[Directory.scala 96:28]
  assign io_read_resp_bits_isDirtyWay = |_isDirtyWay_T; // @[Directory.scala 98:53]
  assign io_read_resp_bits_tagRdVec_0 = ren ? tagArray_io_r_data_0 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_1 = ren ? tagArray_io_r_data_1 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_2 = ren ? tagArray_io_r_data_2 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_3 = ren ? tagArray_io_r_data_3 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_4 = ren ? tagArray_io_r_data_4 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_5 = ren ? tagArray_io_r_data_5 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_6 = ren ? tagArray_io_r_data_6 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_read_resp_bits_tagRdVec_7 = ren ? tagArray_io_r_data_7 : 20'h0; // @[SRAM_1.scala 102:22 103:19 101:32]
  assign io_write_req_ready = 1'h1; // @[Directory.scala 76:29]
  assign tagArray_clock = clock;
  assign tagArray_reset = reset;
  assign tagArray_io_r_addr = rSet; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign tagArray_io_w_en = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  assign tagArray_io_w_addr = wSet; // @[Directory.scala 112:15 SRAM_1.scala 237:19]
  assign tagArray_io_w_data_0 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_1 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_2 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_3 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_4 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_5 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_6 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_data_7 = wTag; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign tagArray_io_w_maskOH = io_write_req_bits_way; // @[Directory.scala 112:15 SRAM_1.scala 239:21]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r_addr = rSet; // @[SRAM_1.scala 102:22 244:{19,19}]
  assign metaArray_io_w_en = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  assign metaArray_io_w_addr = wSet; // @[Directory.scala 112:15 SRAM_1.scala 237:19]
  assign metaArray_io_w_data_0 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_1 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_2 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_3 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_4 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_5 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_6 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_data_7 = io_write_req_bits_meta; // @[Directory.scala 112:15 SRAM_1.scala 238:35]
  assign metaArray_io_w_maskOH = io_write_req_bits_way; // @[Directory.scala 112:15 SRAM_1.scala 239:21]
  assign replaceWay_lfsr_prng_clock = clock;
  assign replaceWay_lfsr_prng_reset = reset;
  always @(posedge clock) begin
    if (_replaceWayReg_T) begin // @[Reg.scala 20:18]
      replaceWayReg <= replaceWay; // @[Reg.scala 20:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_20 < 4'h2)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Error directory write way has multiple valid bit! ==>%d\n    at Directory.scala:69 assert(PopCount(wWay) < 2.U, cf\"Error directory write way has multiple valid bit! ==>${PopCount(wWay)}\")\n"
            ,_T_20); // @[Directory.scala 69:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_20 < 4'h2) & ~reset) begin
          $fatal; // @[Directory.scala 69:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_46 & ~(_T_85 == 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Error chosenWay has multiple valid bit!\n    at Directory.scala:101 assert(PopCount(choseWayOH) === 1.U, \"Error chosenWay has multiple valid bit!\")\n"
            ); // @[Directory.scala 101:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_85 == 4'h1) & _T_46) begin
          $fatal; // @[Directory.scala 101:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wen & _T_46 & ~(_T_20 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: write error, tring to write multiple ways\n    at SRAM_1.scala:235 assert(PopCount(mask) <= 1.U, \"write error, tring to write multiple ways\")\n"
            ); // @[SRAM_1.scala 235:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_20 <= 4'h1) & (wen & _T_46)) begin
          $fatal; // @[SRAM_1.scala 235:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wen & _T_46 & ~(_T_20 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: write error, tring to write multiple ways\n    at SRAM_1.scala:235 assert(PopCount(mask) <= 1.U, \"write error, tring to write multiple ways\")\n"
            ); // @[SRAM_1.scala 235:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_20 <= 4'h1) & (wen & _T_46)) begin
          $fatal; // @[SRAM_1.scala 235:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  replaceWayReg = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input         io_in_0_bits_dirInfo_hit,
  input  [7:0]  io_in_0_bits_dirInfo_chosenWay,
  input         io_in_0_bits_dirInfo_isDirtyWay,
  input  [19:0] io_in_0_bits_dirtyTag,
  input  [31:0] io_in_0_bits_data_0,
  input  [31:0] io_in_0_bits_data_1,
  input  [31:0] io_in_0_bits_data_2,
  input  [31:0] io_in_0_bits_data_3,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input         io_in_1_bits_dirInfo_hit,
  input  [7:0]  io_in_1_bits_dirInfo_chosenWay,
  input         io_in_1_bits_dirInfo_isDirtyWay,
  input  [19:0] io_in_1_bits_dirtyTag,
  input  [31:0] io_in_1_bits_data_0,
  input  [31:0] io_in_1_bits_data_1,
  input  [31:0] io_in_1_bits_data_2,
  input  [31:0] io_in_1_bits_data_3,
  input  [31:0] io_in_1_bits_storeData,
  input  [3:0]  io_in_1_bits_storeMask,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output        io_out_bits_dirInfo_hit,
  output [7:0]  io_out_bits_dirInfo_chosenWay,
  output        io_out_bits_dirInfo_isDirtyWay,
  output [19:0] io_out_bits_dirtyTag,
  output [31:0] io_out_bits_data_0,
  output [31:0] io_out_bits_data_1,
  output [31:0] io_out_bits_data_2,
  output [31:0] io_out_bits_data_3,
  output        io_out_bits_isStore,
  output [31:0] io_out_bits_storeData,
  output [3:0]  io_out_bits_storeMask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_dirInfo_hit = io_in_0_valid ? io_in_0_bits_dirInfo_hit : io_in_1_bits_dirInfo_hit; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_dirInfo_chosenWay = io_in_0_valid ? io_in_0_bits_dirInfo_chosenWay : io_in_1_bits_dirInfo_chosenWay
    ; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_dirInfo_isDirtyWay = io_in_0_valid ? io_in_0_bits_dirInfo_isDirtyWay :
    io_in_1_bits_dirInfo_isDirtyWay; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_dirtyTag = io_in_0_valid ? io_in_0_bits_dirtyTag : io_in_1_bits_dirtyTag; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data_0 = io_in_0_valid ? io_in_0_bits_data_0 : io_in_1_bits_data_0; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data_1 = io_in_0_valid ? io_in_0_bits_data_1 : io_in_1_bits_data_1; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data_2 = io_in_0_valid ? io_in_0_bits_data_2 : io_in_1_bits_data_2; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data_3 = io_in_0_valid ? io_in_0_bits_data_3 : io_in_1_bits_data_3; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_isStore = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_storeData = io_in_0_valid ? 32'h0 : io_in_1_bits_storeData; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_storeMask = io_in_0_valid ? 4'h0 : io_in_1_bits_storeMask; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_1(
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [31:0]  io_in_0_bits_address,
  input  [127:0] io_in_0_bits_data,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [31:0]  io_in_1_bits_address,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_opcode,
  output [31:0]  io_out_bits_address,
  output [127:0] io_out_bits_data
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_opcode = io_in_0_valid ? 3'h2 : 3'h4; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_address = io_in_0_valid ? io_in_0_bits_address : io_in_1_bits_address; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : 128'h0; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_2(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_data,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_data,
  output        io_out_valid,
  output [31:0] io_out_bits_data
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_3(
  input   io_in_0_valid,
  output  io_in_1_ready,
  input   io_in_1_valid,
  output  io_out_valid
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
endmodule
module Arbiter_4(
  input        io_in_0_valid,
  input  [7:0] io_in_0_bits_set,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [7:0] io_in_1_bits_set,
  output       io_out_valid,
  output [7:0] io_out_bits_set
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_set = io_in_0_valid ? io_in_0_bits_set : io_in_1_bits_set; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_5(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  output        io_out_valid,
  output [31:0] io_out_bits_addr
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Arbiter_6(
  input         io_in_0_valid,
  input  [7:0]  io_in_0_bits_set,
  input  [31:0] io_in_0_bits_data_0,
  input  [31:0] io_in_0_bits_data_1,
  input  [31:0] io_in_0_bits_data_2,
  input  [31:0] io_in_0_bits_data_3,
  input  [3:0]  io_in_0_bits_blockMask,
  input  [7:0]  io_in_0_bits_way,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [7:0]  io_in_1_bits_set,
  input  [31:0] io_in_1_bits_data_0,
  input  [31:0] io_in_1_bits_data_1,
  input  [31:0] io_in_1_bits_data_2,
  input  [31:0] io_in_1_bits_data_3,
  input  [7:0]  io_in_1_bits_way,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [7:0]  io_in_2_bits_set,
  input  [31:0] io_in_2_bits_data_0,
  input  [31:0] io_in_2_bits_data_1,
  input  [31:0] io_in_2_bits_data_2,
  input  [31:0] io_in_2_bits_data_3,
  input  [3:0]  io_in_2_bits_blockMask,
  input  [7:0]  io_in_2_bits_way,
  output        io_out_valid,
  output [7:0]  io_out_bits_set,
  output [31:0] io_out_bits_data_0,
  output [31:0] io_out_bits_data_1,
  output [31:0] io_out_bits_data_2,
  output [31:0] io_out_bits_data_3,
  output [3:0]  io_out_bits_blockMask,
  output [7:0]  io_out_bits_way
);
  wire [7:0] _GEN_1 = io_in_1_valid ? io_in_1_bits_set : io_in_2_bits_set; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [31:0] _GEN_3 = io_in_1_valid ? io_in_1_bits_data_0 : io_in_2_bits_data_0; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [31:0] _GEN_4 = io_in_1_valid ? io_in_1_bits_data_1 : io_in_2_bits_data_1; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [31:0] _GEN_5 = io_in_1_valid ? io_in_1_bits_data_2 : io_in_2_bits_data_2; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [31:0] _GEN_6 = io_in_1_valid ? io_in_1_bits_data_3 : io_in_2_bits_data_3; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [3:0] _GEN_7 = io_in_1_valid ? 4'hf : io_in_2_bits_blockMask; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [7:0] _GEN_8 = io_in_1_valid ? io_in_1_bits_way : io_in_2_bits_way; // @[Arbiter.scala 136:15 138:26 140:19]
  wire  grant_2 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_2_ready = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_2 | io_in_2_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_set = io_in_0_valid ? io_in_0_bits_set : _GEN_1; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_data_0 = io_in_0_valid ? io_in_0_bits_data_0 : _GEN_3; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_data_1 = io_in_0_valid ? io_in_0_bits_data_1 : _GEN_4; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_data_2 = io_in_0_valid ? io_in_0_bits_data_2 : _GEN_5; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_data_3 = io_in_0_valid ? io_in_0_bits_data_3 : _GEN_6; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_blockMask = io_in_0_valid ? io_in_0_bits_blockMask : _GEN_7; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_way = io_in_0_valid ? io_in_0_bits_way : _GEN_8; // @[Arbiter.scala 138:26 140:19]
endmodule
module Arbiter_7(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [7:0]  io_in_0_bits_way,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [7:0]  io_in_1_bits_way,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input  [7:0]  io_in_2_bits_way,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [7:0]  io_out_bits_way,
  output [1:0]  io_out_bits_meta
);
  wire [31:0] _GEN_1 = io_in_1_valid ? io_in_1_bits_addr : io_in_2_bits_addr; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [7:0] _GEN_2 = io_in_1_valid ? io_in_1_bits_way : io_in_2_bits_way; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [1:0] _GEN_3 = io_in_1_valid ? 2'h1 : 2'h3; // @[Arbiter.scala 136:15 138:26 140:19]
  wire  grant_2 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_2_ready = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_2 | io_in_2_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_1; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_way = io_in_0_valid ? io_in_0_bits_way : _GEN_2; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_meta = io_in_0_valid ? 2'h3 : _GEN_3; // @[Arbiter.scala 138:26 140:19]
endmodule
module DCache(
  input          clock,
  input          reset,
  output         io_read_req_ready,
  input          io_read_req_valid,
  input  [31:0]  io_read_req_bits_addr,
  output         io_read_resp_valid,
  output [31:0]  io_read_resp_bits_data,
  output         io_write_req_ready,
  input          io_write_req_valid,
  input  [31:0]  io_write_req_bits_addr,
  input  [31:0]  io_write_req_bits_data,
  input  [3:0]   io_write_req_bits_mask,
  output         io_write_resp_valid,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [2:0]   io_tlbus_req_bits_opcode,
  output [31:0]  io_tlbus_req_bits_address,
  output [127:0] io_tlbus_req_bits_data,
  output         io_tlbus_resp_ready,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  loadPipe_clock; // @[DCache.scala 81:26]
  wire  loadPipe_reset; // @[DCache.scala 81:26]
  wire  loadPipe_io_load_req_ready; // @[DCache.scala 81:26]
  wire  loadPipe_io_load_req_valid; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_load_req_bits_addr; // @[DCache.scala 81:26]
  wire  loadPipe_io_load_resp_valid; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_load_resp_bits_data; // @[DCache.scala 81:26]
  wire  loadPipe_io_dir_req_ready; // @[DCache.scala 81:26]
  wire  loadPipe_io_dir_req_valid; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dir_req_bits_addr; // @[DCache.scala 81:26]
  wire  loadPipe_io_dir_resp_bits_hit; // @[DCache.scala 81:26]
  wire [7:0] loadPipe_io_dir_resp_bits_chosenWay; // @[DCache.scala 81:26]
  wire  loadPipe_io_dir_resp_bits_isDirtyWay; // @[DCache.scala 81:26]
  wire [19:0] loadPipe_io_dir_resp_bits_tagRdVec_0; // @[DCache.scala 81:26]
  wire [19:0] loadPipe_io_dir_resp_bits_tagRdVec_1; // @[DCache.scala 81:26]
  wire [19:0] loadPipe_io_dir_resp_bits_tagRdVec_2; // @[DCache.scala 81:26]
  wire [19:0] loadPipe_io_dir_resp_bits_tagRdVec_3; // @[DCache.scala 81:26]
  wire [19:0] loadPipe_io_dir_resp_bits_tagRdVec_4; // @[DCache.scala 81:26]
  wire [19:0] loadPipe_io_dir_resp_bits_tagRdVec_5; // @[DCache.scala 81:26]
  wire [19:0] loadPipe_io_dir_resp_bits_tagRdVec_6; // @[DCache.scala 81:26]
  wire [19:0] loadPipe_io_dir_resp_bits_tagRdVec_7; // @[DCache.scala 81:26]
  wire  loadPipe_io_dataBank_req_ready; // @[DCache.scala 81:26]
  wire  loadPipe_io_dataBank_req_valid; // @[DCache.scala 81:26]
  wire [7:0] loadPipe_io_dataBank_req_bits_set; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_0_0; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_0_1; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_0_2; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_0_3; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_1_0; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_1_1; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_1_2; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_1_3; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_2_0; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_2_1; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_2_2; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_2_3; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_3_0; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_3_1; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_3_2; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_3_3; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_4_0; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_4_1; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_4_2; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_4_3; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_5_0; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_5_1; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_5_2; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_5_3; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_6_0; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_6_1; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_6_2; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_6_3; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_7_0; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_7_1; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_7_2; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_dataBank_resp_7_3; // @[DCache.scala 81:26]
  wire  loadPipe_io_mshr_ready; // @[DCache.scala 81:26]
  wire  loadPipe_io_mshr_valid; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_mshr_bits_addr; // @[DCache.scala 81:26]
  wire  loadPipe_io_mshr_bits_dirInfo_hit; // @[DCache.scala 81:26]
  wire [7:0] loadPipe_io_mshr_bits_dirInfo_chosenWay; // @[DCache.scala 81:26]
  wire  loadPipe_io_mshr_bits_dirInfo_isDirtyWay; // @[DCache.scala 81:26]
  wire [19:0] loadPipe_io_mshr_bits_dirtyTag; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_mshr_bits_data_0; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_mshr_bits_data_1; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_mshr_bits_data_2; // @[DCache.scala 81:26]
  wire [31:0] loadPipe_io_mshr_bits_data_3; // @[DCache.scala 81:26]
  wire  storePipe_clock; // @[DCache.scala 82:27]
  wire  storePipe_reset; // @[DCache.scala 82:27]
  wire  storePipe_io_store_req_ready; // @[DCache.scala 82:27]
  wire  storePipe_io_store_req_valid; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_store_req_bits_addr; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_store_req_bits_data; // @[DCache.scala 82:27]
  wire [3:0] storePipe_io_store_req_bits_mask; // @[DCache.scala 82:27]
  wire  storePipe_io_store_resp_valid; // @[DCache.scala 82:27]
  wire  storePipe_io_dir_read_req_valid; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dir_read_req_bits_addr; // @[DCache.scala 82:27]
  wire  storePipe_io_dir_read_resp_bits_hit; // @[DCache.scala 82:27]
  wire [7:0] storePipe_io_dir_read_resp_bits_chosenWay; // @[DCache.scala 82:27]
  wire  storePipe_io_dir_read_resp_bits_isDirtyWay; // @[DCache.scala 82:27]
  wire [19:0] storePipe_io_dir_read_resp_bits_tagRdVec_0; // @[DCache.scala 82:27]
  wire [19:0] storePipe_io_dir_read_resp_bits_tagRdVec_1; // @[DCache.scala 82:27]
  wire [19:0] storePipe_io_dir_read_resp_bits_tagRdVec_2; // @[DCache.scala 82:27]
  wire [19:0] storePipe_io_dir_read_resp_bits_tagRdVec_3; // @[DCache.scala 82:27]
  wire [19:0] storePipe_io_dir_read_resp_bits_tagRdVec_4; // @[DCache.scala 82:27]
  wire [19:0] storePipe_io_dir_read_resp_bits_tagRdVec_5; // @[DCache.scala 82:27]
  wire [19:0] storePipe_io_dir_read_resp_bits_tagRdVec_6; // @[DCache.scala 82:27]
  wire [19:0] storePipe_io_dir_read_resp_bits_tagRdVec_7; // @[DCache.scala 82:27]
  wire  storePipe_io_dir_write_req_valid; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dir_write_req_bits_addr; // @[DCache.scala 82:27]
  wire [7:0] storePipe_io_dir_write_req_bits_way; // @[DCache.scala 82:27]
  wire  storePipe_io_dataBank_read_req_valid; // @[DCache.scala 82:27]
  wire [7:0] storePipe_io_dataBank_read_req_bits_set; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_0_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_0_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_0_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_0_3; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_1_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_1_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_1_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_1_3; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_2_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_2_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_2_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_2_3; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_3_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_3_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_3_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_3_3; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_4_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_4_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_4_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_4_3; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_5_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_5_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_5_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_5_3; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_6_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_6_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_6_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_6_3; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_7_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_7_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_7_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_read_resp_7_3; // @[DCache.scala 82:27]
  wire  storePipe_io_dataBank_write_req_valid; // @[DCache.scala 82:27]
  wire [7:0] storePipe_io_dataBank_write_req_bits_set; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_write_req_bits_data_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_write_req_bits_data_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_write_req_bits_data_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_dataBank_write_req_bits_data_3; // @[DCache.scala 82:27]
  wire [3:0] storePipe_io_dataBank_write_req_bits_blockMask; // @[DCache.scala 82:27]
  wire [7:0] storePipe_io_dataBank_write_req_bits_way; // @[DCache.scala 82:27]
  wire  storePipe_io_mshr_ready; // @[DCache.scala 82:27]
  wire  storePipe_io_mshr_valid; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_mshr_bits_addr; // @[DCache.scala 82:27]
  wire  storePipe_io_mshr_bits_dirInfo_hit; // @[DCache.scala 82:27]
  wire [7:0] storePipe_io_mshr_bits_dirInfo_chosenWay; // @[DCache.scala 82:27]
  wire  storePipe_io_mshr_bits_dirInfo_isDirtyWay; // @[DCache.scala 82:27]
  wire [19:0] storePipe_io_mshr_bits_dirtyTag; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_mshr_bits_data_0; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_mshr_bits_data_1; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_mshr_bits_data_2; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_mshr_bits_data_3; // @[DCache.scala 82:27]
  wire [31:0] storePipe_io_mshr_bits_storeData; // @[DCache.scala 82:27]
  wire [3:0] storePipe_io_mshr_bits_storeMask; // @[DCache.scala 82:27]
  wire  mshr_clock; // @[DCache.scala 83:22]
  wire  mshr_reset; // @[DCache.scala 83:22]
  wire  mshr_io_req_ready; // @[DCache.scala 83:22]
  wire  mshr_io_req_valid; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_req_bits_addr; // @[DCache.scala 83:22]
  wire  mshr_io_req_bits_dirInfo_hit; // @[DCache.scala 83:22]
  wire [7:0] mshr_io_req_bits_dirInfo_chosenWay; // @[DCache.scala 83:22]
  wire  mshr_io_req_bits_dirInfo_isDirtyWay; // @[DCache.scala 83:22]
  wire [19:0] mshr_io_req_bits_dirtyTag; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_req_bits_data_0; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_req_bits_data_1; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_req_bits_data_2; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_req_bits_data_3; // @[DCache.scala 83:22]
  wire  mshr_io_req_bits_isStore; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_req_bits_storeData; // @[DCache.scala 83:22]
  wire [3:0] mshr_io_req_bits_storeMask; // @[DCache.scala 83:22]
  wire  mshr_io_resp_load_ready; // @[DCache.scala 83:22]
  wire  mshr_io_resp_load_valid; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_resp_load_bits_data; // @[DCache.scala 83:22]
  wire  mshr_io_resp_store_ready; // @[DCache.scala 83:22]
  wire  mshr_io_resp_store_valid; // @[DCache.scala 83:22]
  wire  mshr_io_tasks_refill_req_valid; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_tasks_refill_req_bits_addr; // @[DCache.scala 83:22]
  wire [7:0] mshr_io_tasks_refill_req_bits_chosenWay; // @[DCache.scala 83:22]
  wire  mshr_io_tasks_refill_resp_ready; // @[DCache.scala 83:22]
  wire  mshr_io_tasks_refill_resp_valid; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_tasks_refill_resp_bits_data; // @[DCache.scala 83:22]
  wire  mshr_io_tasks_writeback_req_valid; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_addr; // @[DCache.scala 83:22]
  wire [19:0] mshr_io_tasks_writeback_req_bits_dirtyTag; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_data_0; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_data_1; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_data_2; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_tasks_writeback_req_bits_data_3; // @[DCache.scala 83:22]
  wire  mshr_io_tasks_writeback_resp_ready; // @[DCache.scala 83:22]
  wire  mshr_io_tasks_writeback_resp_valid; // @[DCache.scala 83:22]
  wire  mshr_io_dirWrite_req_ready; // @[DCache.scala 83:22]
  wire  mshr_io_dirWrite_req_valid; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_dirWrite_req_bits_addr; // @[DCache.scala 83:22]
  wire [7:0] mshr_io_dirWrite_req_bits_way; // @[DCache.scala 83:22]
  wire  mshr_io_dataWrite_req_ready; // @[DCache.scala 83:22]
  wire  mshr_io_dataWrite_req_valid; // @[DCache.scala 83:22]
  wire [7:0] mshr_io_dataWrite_req_bits_set; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_dataWrite_req_bits_data_0; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_dataWrite_req_bits_data_1; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_dataWrite_req_bits_data_2; // @[DCache.scala 83:22]
  wire [31:0] mshr_io_dataWrite_req_bits_data_3; // @[DCache.scala 83:22]
  wire [3:0] mshr_io_dataWrite_req_bits_blockMask; // @[DCache.scala 83:22]
  wire [7:0] mshr_io_dataWrite_req_bits_way; // @[DCache.scala 83:22]
  wire  refillPipe_clock; // @[DCache.scala 84:28]
  wire  refillPipe_reset; // @[DCache.scala 84:28]
  wire  refillPipe_io_req_ready; // @[DCache.scala 84:28]
  wire  refillPipe_io_req_valid; // @[DCache.scala 84:28]
  wire [31:0] refillPipe_io_req_bits_addr; // @[DCache.scala 84:28]
  wire [7:0] refillPipe_io_req_bits_chosenWay; // @[DCache.scala 84:28]
  wire  refillPipe_io_resp_valid; // @[DCache.scala 84:28]
  wire [31:0] refillPipe_io_resp_bits_data; // @[DCache.scala 84:28]
  wire  refillPipe_io_tlbus_req_ready; // @[DCache.scala 84:28]
  wire  refillPipe_io_tlbus_req_valid; // @[DCache.scala 84:28]
  wire [127:0] refillPipe_io_tlbus_req_bits_size; // @[DCache.scala 84:28]
  wire [31:0] refillPipe_io_tlbus_req_bits_address; // @[DCache.scala 84:28]
  wire  refillPipe_io_tlbus_resp_ready; // @[DCache.scala 84:28]
  wire  refillPipe_io_tlbus_resp_valid; // @[DCache.scala 84:28]
  wire [2:0] refillPipe_io_tlbus_resp_bits_opcode; // @[DCache.scala 84:28]
  wire [127:0] refillPipe_io_tlbus_resp_bits_data; // @[DCache.scala 84:28]
  wire  refillPipe_io_dirWrite_req_ready; // @[DCache.scala 84:28]
  wire  refillPipe_io_dirWrite_req_valid; // @[DCache.scala 84:28]
  wire [31:0] refillPipe_io_dirWrite_req_bits_addr; // @[DCache.scala 84:28]
  wire [7:0] refillPipe_io_dirWrite_req_bits_way; // @[DCache.scala 84:28]
  wire  refillPipe_io_dataWrite_req_ready; // @[DCache.scala 84:28]
  wire  refillPipe_io_dataWrite_req_valid; // @[DCache.scala 84:28]
  wire [7:0] refillPipe_io_dataWrite_req_bits_set; // @[DCache.scala 84:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_0; // @[DCache.scala 84:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_1; // @[DCache.scala 84:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_2; // @[DCache.scala 84:28]
  wire [31:0] refillPipe_io_dataWrite_req_bits_data_3; // @[DCache.scala 84:28]
  wire [7:0] refillPipe_io_dataWrite_req_bits_way; // @[DCache.scala 84:28]
  wire  wb_clock; // @[DCache.scala 85:20]
  wire  wb_reset; // @[DCache.scala 85:20]
  wire  wb_io_req_ready; // @[DCache.scala 85:20]
  wire  wb_io_req_valid; // @[DCache.scala 85:20]
  wire [31:0] wb_io_req_bits_addr; // @[DCache.scala 85:20]
  wire [19:0] wb_io_req_bits_dirtyTag; // @[DCache.scala 85:20]
  wire [31:0] wb_io_req_bits_data_0; // @[DCache.scala 85:20]
  wire [31:0] wb_io_req_bits_data_1; // @[DCache.scala 85:20]
  wire [31:0] wb_io_req_bits_data_2; // @[DCache.scala 85:20]
  wire [31:0] wb_io_req_bits_data_3; // @[DCache.scala 85:20]
  wire  wb_io_resp_valid; // @[DCache.scala 85:20]
  wire  wb_io_tlbus_req_ready; // @[DCache.scala 85:20]
  wire  wb_io_tlbus_req_valid; // @[DCache.scala 85:20]
  wire [31:0] wb_io_tlbus_req_bits_address; // @[DCache.scala 85:20]
  wire [127:0] wb_io_tlbus_req_bits_data; // @[DCache.scala 85:20]
  wire  wb_io_tlbus_resp_ready; // @[DCache.scala 85:20]
  wire  wb_io_tlbus_resp_valid; // @[DCache.scala 85:20]
  wire  db_clock; // @[DCache.scala 86:20]
  wire  db_reset; // @[DCache.scala 86:20]
  wire  db_io_read_req_ready; // @[DCache.scala 86:20]
  wire  db_io_read_req_valid; // @[DCache.scala 86:20]
  wire [7:0] db_io_read_req_bits_set; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_0_0; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_0_1; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_0_2; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_0_3; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_1_0; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_1_1; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_1_2; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_1_3; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_2_0; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_2_1; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_2_2; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_2_3; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_3_0; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_3_1; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_3_2; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_3_3; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_4_0; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_4_1; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_4_2; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_4_3; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_5_0; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_5_1; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_5_2; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_5_3; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_6_0; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_6_1; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_6_2; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_6_3; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_7_0; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_7_1; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_7_2; // @[DCache.scala 86:20]
  wire [31:0] db_io_read_resp_7_3; // @[DCache.scala 86:20]
  wire  db_io_write_req_ready; // @[DCache.scala 86:20]
  wire  db_io_write_req_valid; // @[DCache.scala 86:20]
  wire [7:0] db_io_write_req_bits_set; // @[DCache.scala 86:20]
  wire [31:0] db_io_write_req_bits_data_0; // @[DCache.scala 86:20]
  wire [31:0] db_io_write_req_bits_data_1; // @[DCache.scala 86:20]
  wire [31:0] db_io_write_req_bits_data_2; // @[DCache.scala 86:20]
  wire [31:0] db_io_write_req_bits_data_3; // @[DCache.scala 86:20]
  wire [3:0] db_io_write_req_bits_blockMask; // @[DCache.scala 86:20]
  wire [7:0] db_io_write_req_bits_way; // @[DCache.scala 86:20]
  wire  dir_clock; // @[DCache.scala 87:21]
  wire  dir_reset; // @[DCache.scala 87:21]
  wire  dir_io_read_req_ready; // @[DCache.scala 87:21]
  wire  dir_io_read_req_valid; // @[DCache.scala 87:21]
  wire [31:0] dir_io_read_req_bits_addr; // @[DCache.scala 87:21]
  wire  dir_io_read_resp_bits_hit; // @[DCache.scala 87:21]
  wire [7:0] dir_io_read_resp_bits_chosenWay; // @[DCache.scala 87:21]
  wire  dir_io_read_resp_bits_isDirtyWay; // @[DCache.scala 87:21]
  wire [19:0] dir_io_read_resp_bits_tagRdVec_0; // @[DCache.scala 87:21]
  wire [19:0] dir_io_read_resp_bits_tagRdVec_1; // @[DCache.scala 87:21]
  wire [19:0] dir_io_read_resp_bits_tagRdVec_2; // @[DCache.scala 87:21]
  wire [19:0] dir_io_read_resp_bits_tagRdVec_3; // @[DCache.scala 87:21]
  wire [19:0] dir_io_read_resp_bits_tagRdVec_4; // @[DCache.scala 87:21]
  wire [19:0] dir_io_read_resp_bits_tagRdVec_5; // @[DCache.scala 87:21]
  wire [19:0] dir_io_read_resp_bits_tagRdVec_6; // @[DCache.scala 87:21]
  wire [19:0] dir_io_read_resp_bits_tagRdVec_7; // @[DCache.scala 87:21]
  wire  dir_io_write_req_ready; // @[DCache.scala 87:21]
  wire  dir_io_write_req_valid; // @[DCache.scala 87:21]
  wire [31:0] dir_io_write_req_bits_addr; // @[DCache.scala 87:21]
  wire [7:0] dir_io_write_req_bits_way; // @[DCache.scala 87:21]
  wire [1:0] dir_io_write_req_bits_meta; // @[DCache.scala 87:21]
  wire  mshrReqArb_io_in_0_ready; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_in_0_valid; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_0_bits_addr; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_in_0_bits_dirInfo_hit; // @[DCache.scala 105:28]
  wire [7:0] mshrReqArb_io_in_0_bits_dirInfo_chosenWay; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_in_0_bits_dirInfo_isDirtyWay; // @[DCache.scala 105:28]
  wire [19:0] mshrReqArb_io_in_0_bits_dirtyTag; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_0_bits_data_0; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_0_bits_data_1; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_0_bits_data_2; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_0_bits_data_3; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_in_1_ready; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_in_1_valid; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_1_bits_addr; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_in_1_bits_dirInfo_hit; // @[DCache.scala 105:28]
  wire [7:0] mshrReqArb_io_in_1_bits_dirInfo_chosenWay; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_in_1_bits_dirInfo_isDirtyWay; // @[DCache.scala 105:28]
  wire [19:0] mshrReqArb_io_in_1_bits_dirtyTag; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_1_bits_data_0; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_1_bits_data_1; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_1_bits_data_2; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_1_bits_data_3; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_in_1_bits_storeData; // @[DCache.scala 105:28]
  wire [3:0] mshrReqArb_io_in_1_bits_storeMask; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_out_ready; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_out_valid; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_out_bits_addr; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_out_bits_dirInfo_hit; // @[DCache.scala 105:28]
  wire [7:0] mshrReqArb_io_out_bits_dirInfo_chosenWay; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_out_bits_dirInfo_isDirtyWay; // @[DCache.scala 105:28]
  wire [19:0] mshrReqArb_io_out_bits_dirtyTag; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_out_bits_data_0; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_out_bits_data_1; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_out_bits_data_2; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_out_bits_data_3; // @[DCache.scala 105:28]
  wire  mshrReqArb_io_out_bits_isStore; // @[DCache.scala 105:28]
  wire [31:0] mshrReqArb_io_out_bits_storeData; // @[DCache.scala 105:28]
  wire [3:0] mshrReqArb_io_out_bits_storeMask; // @[DCache.scala 105:28]
  wire  tlbusReqArb_io_in_0_ready; // @[DCache.scala 110:29]
  wire  tlbusReqArb_io_in_0_valid; // @[DCache.scala 110:29]
  wire [31:0] tlbusReqArb_io_in_0_bits_address; // @[DCache.scala 110:29]
  wire [127:0] tlbusReqArb_io_in_0_bits_data; // @[DCache.scala 110:29]
  wire  tlbusReqArb_io_in_1_ready; // @[DCache.scala 110:29]
  wire  tlbusReqArb_io_in_1_valid; // @[DCache.scala 110:29]
  wire [31:0] tlbusReqArb_io_in_1_bits_address; // @[DCache.scala 110:29]
  wire  tlbusReqArb_io_out_ready; // @[DCache.scala 110:29]
  wire  tlbusReqArb_io_out_valid; // @[DCache.scala 110:29]
  wire [2:0] tlbusReqArb_io_out_bits_opcode; // @[DCache.scala 110:29]
  wire [31:0] tlbusReqArb_io_out_bits_address; // @[DCache.scala 110:29]
  wire [127:0] tlbusReqArb_io_out_bits_data; // @[DCache.scala 110:29]
  wire  loadRespArb_io_in_0_valid; // @[DCache.scala 122:29]
  wire [31:0] loadRespArb_io_in_0_bits_data; // @[DCache.scala 122:29]
  wire  loadRespArb_io_in_1_ready; // @[DCache.scala 122:29]
  wire  loadRespArb_io_in_1_valid; // @[DCache.scala 122:29]
  wire [31:0] loadRespArb_io_in_1_bits_data; // @[DCache.scala 122:29]
  wire  loadRespArb_io_out_valid; // @[DCache.scala 122:29]
  wire [31:0] loadRespArb_io_out_bits_data; // @[DCache.scala 122:29]
  wire  storeRespArb_io_in_0_valid; // @[DCache.scala 127:30]
  wire  storeRespArb_io_in_1_ready; // @[DCache.scala 127:30]
  wire  storeRespArb_io_in_1_valid; // @[DCache.scala 127:30]
  wire  storeRespArb_io_out_valid; // @[DCache.scala 127:30]
  wire  dbRdReqArb_io_in_0_valid; // @[DCache.scala 133:28]
  wire [7:0] dbRdReqArb_io_in_0_bits_set; // @[DCache.scala 133:28]
  wire  dbRdReqArb_io_in_1_ready; // @[DCache.scala 133:28]
  wire  dbRdReqArb_io_in_1_valid; // @[DCache.scala 133:28]
  wire [7:0] dbRdReqArb_io_in_1_bits_set; // @[DCache.scala 133:28]
  wire  dbRdReqArb_io_out_valid; // @[DCache.scala 133:28]
  wire [7:0] dbRdReqArb_io_out_bits_set; // @[DCache.scala 133:28]
  wire  dirRdReqArb_io_in_0_valid; // @[DCache.scala 138:29]
  wire [31:0] dirRdReqArb_io_in_0_bits_addr; // @[DCache.scala 138:29]
  wire  dirRdReqArb_io_in_1_ready; // @[DCache.scala 138:29]
  wire  dirRdReqArb_io_in_1_valid; // @[DCache.scala 138:29]
  wire [31:0] dirRdReqArb_io_in_1_bits_addr; // @[DCache.scala 138:29]
  wire  dirRdReqArb_io_out_valid; // @[DCache.scala 138:29]
  wire [31:0] dirRdReqArb_io_out_bits_addr; // @[DCache.scala 138:29]
  wire  dataBankWrArb_io_in_0_valid; // @[DCache.scala 144:31]
  wire [7:0] dataBankWrArb_io_in_0_bits_set; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_0_bits_data_0; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_0_bits_data_1; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_0_bits_data_2; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_0_bits_data_3; // @[DCache.scala 144:31]
  wire [3:0] dataBankWrArb_io_in_0_bits_blockMask; // @[DCache.scala 144:31]
  wire [7:0] dataBankWrArb_io_in_0_bits_way; // @[DCache.scala 144:31]
  wire  dataBankWrArb_io_in_1_ready; // @[DCache.scala 144:31]
  wire  dataBankWrArb_io_in_1_valid; // @[DCache.scala 144:31]
  wire [7:0] dataBankWrArb_io_in_1_bits_set; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_1_bits_data_0; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_1_bits_data_1; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_1_bits_data_2; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_1_bits_data_3; // @[DCache.scala 144:31]
  wire [7:0] dataBankWrArb_io_in_1_bits_way; // @[DCache.scala 144:31]
  wire  dataBankWrArb_io_in_2_ready; // @[DCache.scala 144:31]
  wire  dataBankWrArb_io_in_2_valid; // @[DCache.scala 144:31]
  wire [7:0] dataBankWrArb_io_in_2_bits_set; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_2_bits_data_0; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_2_bits_data_1; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_2_bits_data_2; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_in_2_bits_data_3; // @[DCache.scala 144:31]
  wire [3:0] dataBankWrArb_io_in_2_bits_blockMask; // @[DCache.scala 144:31]
  wire [7:0] dataBankWrArb_io_in_2_bits_way; // @[DCache.scala 144:31]
  wire  dataBankWrArb_io_out_valid; // @[DCache.scala 144:31]
  wire [7:0] dataBankWrArb_io_out_bits_set; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_out_bits_data_0; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_out_bits_data_1; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_out_bits_data_2; // @[DCache.scala 144:31]
  wire [31:0] dataBankWrArb_io_out_bits_data_3; // @[DCache.scala 144:31]
  wire [3:0] dataBankWrArb_io_out_bits_blockMask; // @[DCache.scala 144:31]
  wire [7:0] dataBankWrArb_io_out_bits_way; // @[DCache.scala 144:31]
  wire  dirWrArb_io_in_0_valid; // @[DCache.scala 150:26]
  wire [31:0] dirWrArb_io_in_0_bits_addr; // @[DCache.scala 150:26]
  wire [7:0] dirWrArb_io_in_0_bits_way; // @[DCache.scala 150:26]
  wire  dirWrArb_io_in_1_ready; // @[DCache.scala 150:26]
  wire  dirWrArb_io_in_1_valid; // @[DCache.scala 150:26]
  wire [31:0] dirWrArb_io_in_1_bits_addr; // @[DCache.scala 150:26]
  wire [7:0] dirWrArb_io_in_1_bits_way; // @[DCache.scala 150:26]
  wire  dirWrArb_io_in_2_ready; // @[DCache.scala 150:26]
  wire  dirWrArb_io_in_2_valid; // @[DCache.scala 150:26]
  wire [31:0] dirWrArb_io_in_2_bits_addr; // @[DCache.scala 150:26]
  wire [7:0] dirWrArb_io_in_2_bits_way; // @[DCache.scala 150:26]
  wire  dirWrArb_io_out_valid; // @[DCache.scala 150:26]
  wire [31:0] dirWrArb_io_out_bits_addr; // @[DCache.scala 150:26]
  wire [7:0] dirWrArb_io_out_bits_way; // @[DCache.scala 150:26]
  wire [1:0] dirWrArb_io_out_bits_meta; // @[DCache.scala 150:26]
  wire  _T = io_read_req_ready & io_read_req_valid; // @[Decoupled.scala 51:35]
  reg [63:0] c; // @[util.scala 162:24]
  wire [63:0] _c_T_1 = c + 64'h1; // @[util.scala 163:16]
  reg [63:0] c_1; // @[util.scala 162:24]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[util.scala 163:16]
  wire  _T_6 = io_write_req_ready & io_write_req_valid; // @[Decoupled.scala 51:35]
  reg [63:0] c_2; // @[util.scala 162:24]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[util.scala 163:16]
  reg [63:0] c_3; // @[util.scala 162:24]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[util.scala 163:16]
  wire  _T_12 = io_tlbus_req_ready & io_tlbus_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_14 = _T_12 & io_tlbus_req_bits_opcode == 3'h2; // @[DCache.scala 162:54]
  reg [63:0] c_4; // @[util.scala 162:24]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[util.scala 163:16]
  wire  _T_17 = io_tlbus_resp_ready & io_tlbus_resp_valid; // @[Decoupled.scala 51:35]
  wire  _T_19 = _T_17 & io_tlbus_resp_bits_opcode == 3'h1; // @[DCache.scala 163:55]
  reg [63:0] c_5; // @[util.scala 162:24]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[util.scala 163:16]
  LoadPipe loadPipe ( // @[DCache.scala 81:26]
    .clock(loadPipe_clock),
    .reset(loadPipe_reset),
    .io_load_req_ready(loadPipe_io_load_req_ready),
    .io_load_req_valid(loadPipe_io_load_req_valid),
    .io_load_req_bits_addr(loadPipe_io_load_req_bits_addr),
    .io_load_resp_valid(loadPipe_io_load_resp_valid),
    .io_load_resp_bits_data(loadPipe_io_load_resp_bits_data),
    .io_dir_req_ready(loadPipe_io_dir_req_ready),
    .io_dir_req_valid(loadPipe_io_dir_req_valid),
    .io_dir_req_bits_addr(loadPipe_io_dir_req_bits_addr),
    .io_dir_resp_bits_hit(loadPipe_io_dir_resp_bits_hit),
    .io_dir_resp_bits_chosenWay(loadPipe_io_dir_resp_bits_chosenWay),
    .io_dir_resp_bits_isDirtyWay(loadPipe_io_dir_resp_bits_isDirtyWay),
    .io_dir_resp_bits_tagRdVec_0(loadPipe_io_dir_resp_bits_tagRdVec_0),
    .io_dir_resp_bits_tagRdVec_1(loadPipe_io_dir_resp_bits_tagRdVec_1),
    .io_dir_resp_bits_tagRdVec_2(loadPipe_io_dir_resp_bits_tagRdVec_2),
    .io_dir_resp_bits_tagRdVec_3(loadPipe_io_dir_resp_bits_tagRdVec_3),
    .io_dir_resp_bits_tagRdVec_4(loadPipe_io_dir_resp_bits_tagRdVec_4),
    .io_dir_resp_bits_tagRdVec_5(loadPipe_io_dir_resp_bits_tagRdVec_5),
    .io_dir_resp_bits_tagRdVec_6(loadPipe_io_dir_resp_bits_tagRdVec_6),
    .io_dir_resp_bits_tagRdVec_7(loadPipe_io_dir_resp_bits_tagRdVec_7),
    .io_dataBank_req_ready(loadPipe_io_dataBank_req_ready),
    .io_dataBank_req_valid(loadPipe_io_dataBank_req_valid),
    .io_dataBank_req_bits_set(loadPipe_io_dataBank_req_bits_set),
    .io_dataBank_resp_0_0(loadPipe_io_dataBank_resp_0_0),
    .io_dataBank_resp_0_1(loadPipe_io_dataBank_resp_0_1),
    .io_dataBank_resp_0_2(loadPipe_io_dataBank_resp_0_2),
    .io_dataBank_resp_0_3(loadPipe_io_dataBank_resp_0_3),
    .io_dataBank_resp_1_0(loadPipe_io_dataBank_resp_1_0),
    .io_dataBank_resp_1_1(loadPipe_io_dataBank_resp_1_1),
    .io_dataBank_resp_1_2(loadPipe_io_dataBank_resp_1_2),
    .io_dataBank_resp_1_3(loadPipe_io_dataBank_resp_1_3),
    .io_dataBank_resp_2_0(loadPipe_io_dataBank_resp_2_0),
    .io_dataBank_resp_2_1(loadPipe_io_dataBank_resp_2_1),
    .io_dataBank_resp_2_2(loadPipe_io_dataBank_resp_2_2),
    .io_dataBank_resp_2_3(loadPipe_io_dataBank_resp_2_3),
    .io_dataBank_resp_3_0(loadPipe_io_dataBank_resp_3_0),
    .io_dataBank_resp_3_1(loadPipe_io_dataBank_resp_3_1),
    .io_dataBank_resp_3_2(loadPipe_io_dataBank_resp_3_2),
    .io_dataBank_resp_3_3(loadPipe_io_dataBank_resp_3_3),
    .io_dataBank_resp_4_0(loadPipe_io_dataBank_resp_4_0),
    .io_dataBank_resp_4_1(loadPipe_io_dataBank_resp_4_1),
    .io_dataBank_resp_4_2(loadPipe_io_dataBank_resp_4_2),
    .io_dataBank_resp_4_3(loadPipe_io_dataBank_resp_4_3),
    .io_dataBank_resp_5_0(loadPipe_io_dataBank_resp_5_0),
    .io_dataBank_resp_5_1(loadPipe_io_dataBank_resp_5_1),
    .io_dataBank_resp_5_2(loadPipe_io_dataBank_resp_5_2),
    .io_dataBank_resp_5_3(loadPipe_io_dataBank_resp_5_3),
    .io_dataBank_resp_6_0(loadPipe_io_dataBank_resp_6_0),
    .io_dataBank_resp_6_1(loadPipe_io_dataBank_resp_6_1),
    .io_dataBank_resp_6_2(loadPipe_io_dataBank_resp_6_2),
    .io_dataBank_resp_6_3(loadPipe_io_dataBank_resp_6_3),
    .io_dataBank_resp_7_0(loadPipe_io_dataBank_resp_7_0),
    .io_dataBank_resp_7_1(loadPipe_io_dataBank_resp_7_1),
    .io_dataBank_resp_7_2(loadPipe_io_dataBank_resp_7_2),
    .io_dataBank_resp_7_3(loadPipe_io_dataBank_resp_7_3),
    .io_mshr_ready(loadPipe_io_mshr_ready),
    .io_mshr_valid(loadPipe_io_mshr_valid),
    .io_mshr_bits_addr(loadPipe_io_mshr_bits_addr),
    .io_mshr_bits_dirInfo_hit(loadPipe_io_mshr_bits_dirInfo_hit),
    .io_mshr_bits_dirInfo_chosenWay(loadPipe_io_mshr_bits_dirInfo_chosenWay),
    .io_mshr_bits_dirInfo_isDirtyWay(loadPipe_io_mshr_bits_dirInfo_isDirtyWay),
    .io_mshr_bits_dirtyTag(loadPipe_io_mshr_bits_dirtyTag),
    .io_mshr_bits_data_0(loadPipe_io_mshr_bits_data_0),
    .io_mshr_bits_data_1(loadPipe_io_mshr_bits_data_1),
    .io_mshr_bits_data_2(loadPipe_io_mshr_bits_data_2),
    .io_mshr_bits_data_3(loadPipe_io_mshr_bits_data_3)
  );
  StorePipe storePipe ( // @[DCache.scala 82:27]
    .clock(storePipe_clock),
    .reset(storePipe_reset),
    .io_store_req_ready(storePipe_io_store_req_ready),
    .io_store_req_valid(storePipe_io_store_req_valid),
    .io_store_req_bits_addr(storePipe_io_store_req_bits_addr),
    .io_store_req_bits_data(storePipe_io_store_req_bits_data),
    .io_store_req_bits_mask(storePipe_io_store_req_bits_mask),
    .io_store_resp_valid(storePipe_io_store_resp_valid),
    .io_dir_read_req_valid(storePipe_io_dir_read_req_valid),
    .io_dir_read_req_bits_addr(storePipe_io_dir_read_req_bits_addr),
    .io_dir_read_resp_bits_hit(storePipe_io_dir_read_resp_bits_hit),
    .io_dir_read_resp_bits_chosenWay(storePipe_io_dir_read_resp_bits_chosenWay),
    .io_dir_read_resp_bits_isDirtyWay(storePipe_io_dir_read_resp_bits_isDirtyWay),
    .io_dir_read_resp_bits_tagRdVec_0(storePipe_io_dir_read_resp_bits_tagRdVec_0),
    .io_dir_read_resp_bits_tagRdVec_1(storePipe_io_dir_read_resp_bits_tagRdVec_1),
    .io_dir_read_resp_bits_tagRdVec_2(storePipe_io_dir_read_resp_bits_tagRdVec_2),
    .io_dir_read_resp_bits_tagRdVec_3(storePipe_io_dir_read_resp_bits_tagRdVec_3),
    .io_dir_read_resp_bits_tagRdVec_4(storePipe_io_dir_read_resp_bits_tagRdVec_4),
    .io_dir_read_resp_bits_tagRdVec_5(storePipe_io_dir_read_resp_bits_tagRdVec_5),
    .io_dir_read_resp_bits_tagRdVec_6(storePipe_io_dir_read_resp_bits_tagRdVec_6),
    .io_dir_read_resp_bits_tagRdVec_7(storePipe_io_dir_read_resp_bits_tagRdVec_7),
    .io_dir_write_req_valid(storePipe_io_dir_write_req_valid),
    .io_dir_write_req_bits_addr(storePipe_io_dir_write_req_bits_addr),
    .io_dir_write_req_bits_way(storePipe_io_dir_write_req_bits_way),
    .io_dataBank_read_req_valid(storePipe_io_dataBank_read_req_valid),
    .io_dataBank_read_req_bits_set(storePipe_io_dataBank_read_req_bits_set),
    .io_dataBank_read_resp_0_0(storePipe_io_dataBank_read_resp_0_0),
    .io_dataBank_read_resp_0_1(storePipe_io_dataBank_read_resp_0_1),
    .io_dataBank_read_resp_0_2(storePipe_io_dataBank_read_resp_0_2),
    .io_dataBank_read_resp_0_3(storePipe_io_dataBank_read_resp_0_3),
    .io_dataBank_read_resp_1_0(storePipe_io_dataBank_read_resp_1_0),
    .io_dataBank_read_resp_1_1(storePipe_io_dataBank_read_resp_1_1),
    .io_dataBank_read_resp_1_2(storePipe_io_dataBank_read_resp_1_2),
    .io_dataBank_read_resp_1_3(storePipe_io_dataBank_read_resp_1_3),
    .io_dataBank_read_resp_2_0(storePipe_io_dataBank_read_resp_2_0),
    .io_dataBank_read_resp_2_1(storePipe_io_dataBank_read_resp_2_1),
    .io_dataBank_read_resp_2_2(storePipe_io_dataBank_read_resp_2_2),
    .io_dataBank_read_resp_2_3(storePipe_io_dataBank_read_resp_2_3),
    .io_dataBank_read_resp_3_0(storePipe_io_dataBank_read_resp_3_0),
    .io_dataBank_read_resp_3_1(storePipe_io_dataBank_read_resp_3_1),
    .io_dataBank_read_resp_3_2(storePipe_io_dataBank_read_resp_3_2),
    .io_dataBank_read_resp_3_3(storePipe_io_dataBank_read_resp_3_3),
    .io_dataBank_read_resp_4_0(storePipe_io_dataBank_read_resp_4_0),
    .io_dataBank_read_resp_4_1(storePipe_io_dataBank_read_resp_4_1),
    .io_dataBank_read_resp_4_2(storePipe_io_dataBank_read_resp_4_2),
    .io_dataBank_read_resp_4_3(storePipe_io_dataBank_read_resp_4_3),
    .io_dataBank_read_resp_5_0(storePipe_io_dataBank_read_resp_5_0),
    .io_dataBank_read_resp_5_1(storePipe_io_dataBank_read_resp_5_1),
    .io_dataBank_read_resp_5_2(storePipe_io_dataBank_read_resp_5_2),
    .io_dataBank_read_resp_5_3(storePipe_io_dataBank_read_resp_5_3),
    .io_dataBank_read_resp_6_0(storePipe_io_dataBank_read_resp_6_0),
    .io_dataBank_read_resp_6_1(storePipe_io_dataBank_read_resp_6_1),
    .io_dataBank_read_resp_6_2(storePipe_io_dataBank_read_resp_6_2),
    .io_dataBank_read_resp_6_3(storePipe_io_dataBank_read_resp_6_3),
    .io_dataBank_read_resp_7_0(storePipe_io_dataBank_read_resp_7_0),
    .io_dataBank_read_resp_7_1(storePipe_io_dataBank_read_resp_7_1),
    .io_dataBank_read_resp_7_2(storePipe_io_dataBank_read_resp_7_2),
    .io_dataBank_read_resp_7_3(storePipe_io_dataBank_read_resp_7_3),
    .io_dataBank_write_req_valid(storePipe_io_dataBank_write_req_valid),
    .io_dataBank_write_req_bits_set(storePipe_io_dataBank_write_req_bits_set),
    .io_dataBank_write_req_bits_data_0(storePipe_io_dataBank_write_req_bits_data_0),
    .io_dataBank_write_req_bits_data_1(storePipe_io_dataBank_write_req_bits_data_1),
    .io_dataBank_write_req_bits_data_2(storePipe_io_dataBank_write_req_bits_data_2),
    .io_dataBank_write_req_bits_data_3(storePipe_io_dataBank_write_req_bits_data_3),
    .io_dataBank_write_req_bits_blockMask(storePipe_io_dataBank_write_req_bits_blockMask),
    .io_dataBank_write_req_bits_way(storePipe_io_dataBank_write_req_bits_way),
    .io_mshr_ready(storePipe_io_mshr_ready),
    .io_mshr_valid(storePipe_io_mshr_valid),
    .io_mshr_bits_addr(storePipe_io_mshr_bits_addr),
    .io_mshr_bits_dirInfo_hit(storePipe_io_mshr_bits_dirInfo_hit),
    .io_mshr_bits_dirInfo_chosenWay(storePipe_io_mshr_bits_dirInfo_chosenWay),
    .io_mshr_bits_dirInfo_isDirtyWay(storePipe_io_mshr_bits_dirInfo_isDirtyWay),
    .io_mshr_bits_dirtyTag(storePipe_io_mshr_bits_dirtyTag),
    .io_mshr_bits_data_0(storePipe_io_mshr_bits_data_0),
    .io_mshr_bits_data_1(storePipe_io_mshr_bits_data_1),
    .io_mshr_bits_data_2(storePipe_io_mshr_bits_data_2),
    .io_mshr_bits_data_3(storePipe_io_mshr_bits_data_3),
    .io_mshr_bits_storeData(storePipe_io_mshr_bits_storeData),
    .io_mshr_bits_storeMask(storePipe_io_mshr_bits_storeMask)
  );
  MSHR mshr ( // @[DCache.scala 83:22]
    .clock(mshr_clock),
    .reset(mshr_reset),
    .io_req_ready(mshr_io_req_ready),
    .io_req_valid(mshr_io_req_valid),
    .io_req_bits_addr(mshr_io_req_bits_addr),
    .io_req_bits_dirInfo_hit(mshr_io_req_bits_dirInfo_hit),
    .io_req_bits_dirInfo_chosenWay(mshr_io_req_bits_dirInfo_chosenWay),
    .io_req_bits_dirInfo_isDirtyWay(mshr_io_req_bits_dirInfo_isDirtyWay),
    .io_req_bits_dirtyTag(mshr_io_req_bits_dirtyTag),
    .io_req_bits_data_0(mshr_io_req_bits_data_0),
    .io_req_bits_data_1(mshr_io_req_bits_data_1),
    .io_req_bits_data_2(mshr_io_req_bits_data_2),
    .io_req_bits_data_3(mshr_io_req_bits_data_3),
    .io_req_bits_isStore(mshr_io_req_bits_isStore),
    .io_req_bits_storeData(mshr_io_req_bits_storeData),
    .io_req_bits_storeMask(mshr_io_req_bits_storeMask),
    .io_resp_load_ready(mshr_io_resp_load_ready),
    .io_resp_load_valid(mshr_io_resp_load_valid),
    .io_resp_load_bits_data(mshr_io_resp_load_bits_data),
    .io_resp_store_ready(mshr_io_resp_store_ready),
    .io_resp_store_valid(mshr_io_resp_store_valid),
    .io_tasks_refill_req_valid(mshr_io_tasks_refill_req_valid),
    .io_tasks_refill_req_bits_addr(mshr_io_tasks_refill_req_bits_addr),
    .io_tasks_refill_req_bits_chosenWay(mshr_io_tasks_refill_req_bits_chosenWay),
    .io_tasks_refill_resp_ready(mshr_io_tasks_refill_resp_ready),
    .io_tasks_refill_resp_valid(mshr_io_tasks_refill_resp_valid),
    .io_tasks_refill_resp_bits_data(mshr_io_tasks_refill_resp_bits_data),
    .io_tasks_writeback_req_valid(mshr_io_tasks_writeback_req_valid),
    .io_tasks_writeback_req_bits_addr(mshr_io_tasks_writeback_req_bits_addr),
    .io_tasks_writeback_req_bits_dirtyTag(mshr_io_tasks_writeback_req_bits_dirtyTag),
    .io_tasks_writeback_req_bits_data_0(mshr_io_tasks_writeback_req_bits_data_0),
    .io_tasks_writeback_req_bits_data_1(mshr_io_tasks_writeback_req_bits_data_1),
    .io_tasks_writeback_req_bits_data_2(mshr_io_tasks_writeback_req_bits_data_2),
    .io_tasks_writeback_req_bits_data_3(mshr_io_tasks_writeback_req_bits_data_3),
    .io_tasks_writeback_resp_ready(mshr_io_tasks_writeback_resp_ready),
    .io_tasks_writeback_resp_valid(mshr_io_tasks_writeback_resp_valid),
    .io_dirWrite_req_ready(mshr_io_dirWrite_req_ready),
    .io_dirWrite_req_valid(mshr_io_dirWrite_req_valid),
    .io_dirWrite_req_bits_addr(mshr_io_dirWrite_req_bits_addr),
    .io_dirWrite_req_bits_way(mshr_io_dirWrite_req_bits_way),
    .io_dataWrite_req_ready(mshr_io_dataWrite_req_ready),
    .io_dataWrite_req_valid(mshr_io_dataWrite_req_valid),
    .io_dataWrite_req_bits_set(mshr_io_dataWrite_req_bits_set),
    .io_dataWrite_req_bits_data_0(mshr_io_dataWrite_req_bits_data_0),
    .io_dataWrite_req_bits_data_1(mshr_io_dataWrite_req_bits_data_1),
    .io_dataWrite_req_bits_data_2(mshr_io_dataWrite_req_bits_data_2),
    .io_dataWrite_req_bits_data_3(mshr_io_dataWrite_req_bits_data_3),
    .io_dataWrite_req_bits_blockMask(mshr_io_dataWrite_req_bits_blockMask),
    .io_dataWrite_req_bits_way(mshr_io_dataWrite_req_bits_way)
  );
  RefillPipe_1 refillPipe ( // @[DCache.scala 84:28]
    .clock(refillPipe_clock),
    .reset(refillPipe_reset),
    .io_req_ready(refillPipe_io_req_ready),
    .io_req_valid(refillPipe_io_req_valid),
    .io_req_bits_addr(refillPipe_io_req_bits_addr),
    .io_req_bits_chosenWay(refillPipe_io_req_bits_chosenWay),
    .io_resp_valid(refillPipe_io_resp_valid),
    .io_resp_bits_data(refillPipe_io_resp_bits_data),
    .io_tlbus_req_ready(refillPipe_io_tlbus_req_ready),
    .io_tlbus_req_valid(refillPipe_io_tlbus_req_valid),
    .io_tlbus_req_bits_size(refillPipe_io_tlbus_req_bits_size),
    .io_tlbus_req_bits_address(refillPipe_io_tlbus_req_bits_address),
    .io_tlbus_resp_ready(refillPipe_io_tlbus_resp_ready),
    .io_tlbus_resp_valid(refillPipe_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(refillPipe_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(refillPipe_io_tlbus_resp_bits_data),
    .io_dirWrite_req_ready(refillPipe_io_dirWrite_req_ready),
    .io_dirWrite_req_valid(refillPipe_io_dirWrite_req_valid),
    .io_dirWrite_req_bits_addr(refillPipe_io_dirWrite_req_bits_addr),
    .io_dirWrite_req_bits_way(refillPipe_io_dirWrite_req_bits_way),
    .io_dataWrite_req_ready(refillPipe_io_dataWrite_req_ready),
    .io_dataWrite_req_valid(refillPipe_io_dataWrite_req_valid),
    .io_dataWrite_req_bits_set(refillPipe_io_dataWrite_req_bits_set),
    .io_dataWrite_req_bits_data_0(refillPipe_io_dataWrite_req_bits_data_0),
    .io_dataWrite_req_bits_data_1(refillPipe_io_dataWrite_req_bits_data_1),
    .io_dataWrite_req_bits_data_2(refillPipe_io_dataWrite_req_bits_data_2),
    .io_dataWrite_req_bits_data_3(refillPipe_io_dataWrite_req_bits_data_3),
    .io_dataWrite_req_bits_way(refillPipe_io_dataWrite_req_bits_way)
  );
  WritebackQueue wb ( // @[DCache.scala 85:20]
    .clock(wb_clock),
    .reset(wb_reset),
    .io_req_ready(wb_io_req_ready),
    .io_req_valid(wb_io_req_valid),
    .io_req_bits_addr(wb_io_req_bits_addr),
    .io_req_bits_dirtyTag(wb_io_req_bits_dirtyTag),
    .io_req_bits_data_0(wb_io_req_bits_data_0),
    .io_req_bits_data_1(wb_io_req_bits_data_1),
    .io_req_bits_data_2(wb_io_req_bits_data_2),
    .io_req_bits_data_3(wb_io_req_bits_data_3),
    .io_resp_valid(wb_io_resp_valid),
    .io_tlbus_req_ready(wb_io_tlbus_req_ready),
    .io_tlbus_req_valid(wb_io_tlbus_req_valid),
    .io_tlbus_req_bits_address(wb_io_tlbus_req_bits_address),
    .io_tlbus_req_bits_data(wb_io_tlbus_req_bits_data),
    .io_tlbus_resp_ready(wb_io_tlbus_resp_ready),
    .io_tlbus_resp_valid(wb_io_tlbus_resp_valid)
  );
  DataBankArray_1 db ( // @[DCache.scala 86:20]
    .clock(db_clock),
    .reset(db_reset),
    .io_read_req_ready(db_io_read_req_ready),
    .io_read_req_valid(db_io_read_req_valid),
    .io_read_req_bits_set(db_io_read_req_bits_set),
    .io_read_resp_0_0(db_io_read_resp_0_0),
    .io_read_resp_0_1(db_io_read_resp_0_1),
    .io_read_resp_0_2(db_io_read_resp_0_2),
    .io_read_resp_0_3(db_io_read_resp_0_3),
    .io_read_resp_1_0(db_io_read_resp_1_0),
    .io_read_resp_1_1(db_io_read_resp_1_1),
    .io_read_resp_1_2(db_io_read_resp_1_2),
    .io_read_resp_1_3(db_io_read_resp_1_3),
    .io_read_resp_2_0(db_io_read_resp_2_0),
    .io_read_resp_2_1(db_io_read_resp_2_1),
    .io_read_resp_2_2(db_io_read_resp_2_2),
    .io_read_resp_2_3(db_io_read_resp_2_3),
    .io_read_resp_3_0(db_io_read_resp_3_0),
    .io_read_resp_3_1(db_io_read_resp_3_1),
    .io_read_resp_3_2(db_io_read_resp_3_2),
    .io_read_resp_3_3(db_io_read_resp_3_3),
    .io_read_resp_4_0(db_io_read_resp_4_0),
    .io_read_resp_4_1(db_io_read_resp_4_1),
    .io_read_resp_4_2(db_io_read_resp_4_2),
    .io_read_resp_4_3(db_io_read_resp_4_3),
    .io_read_resp_5_0(db_io_read_resp_5_0),
    .io_read_resp_5_1(db_io_read_resp_5_1),
    .io_read_resp_5_2(db_io_read_resp_5_2),
    .io_read_resp_5_3(db_io_read_resp_5_3),
    .io_read_resp_6_0(db_io_read_resp_6_0),
    .io_read_resp_6_1(db_io_read_resp_6_1),
    .io_read_resp_6_2(db_io_read_resp_6_2),
    .io_read_resp_6_3(db_io_read_resp_6_3),
    .io_read_resp_7_0(db_io_read_resp_7_0),
    .io_read_resp_7_1(db_io_read_resp_7_1),
    .io_read_resp_7_2(db_io_read_resp_7_2),
    .io_read_resp_7_3(db_io_read_resp_7_3),
    .io_write_req_ready(db_io_write_req_ready),
    .io_write_req_valid(db_io_write_req_valid),
    .io_write_req_bits_set(db_io_write_req_bits_set),
    .io_write_req_bits_data_0(db_io_write_req_bits_data_0),
    .io_write_req_bits_data_1(db_io_write_req_bits_data_1),
    .io_write_req_bits_data_2(db_io_write_req_bits_data_2),
    .io_write_req_bits_data_3(db_io_write_req_bits_data_3),
    .io_write_req_bits_blockMask(db_io_write_req_bits_blockMask),
    .io_write_req_bits_way(db_io_write_req_bits_way)
  );
  DCacheDirectory_1 dir ( // @[DCache.scala 87:21]
    .clock(dir_clock),
    .reset(dir_reset),
    .io_read_req_ready(dir_io_read_req_ready),
    .io_read_req_valid(dir_io_read_req_valid),
    .io_read_req_bits_addr(dir_io_read_req_bits_addr),
    .io_read_resp_bits_hit(dir_io_read_resp_bits_hit),
    .io_read_resp_bits_chosenWay(dir_io_read_resp_bits_chosenWay),
    .io_read_resp_bits_isDirtyWay(dir_io_read_resp_bits_isDirtyWay),
    .io_read_resp_bits_tagRdVec_0(dir_io_read_resp_bits_tagRdVec_0),
    .io_read_resp_bits_tagRdVec_1(dir_io_read_resp_bits_tagRdVec_1),
    .io_read_resp_bits_tagRdVec_2(dir_io_read_resp_bits_tagRdVec_2),
    .io_read_resp_bits_tagRdVec_3(dir_io_read_resp_bits_tagRdVec_3),
    .io_read_resp_bits_tagRdVec_4(dir_io_read_resp_bits_tagRdVec_4),
    .io_read_resp_bits_tagRdVec_5(dir_io_read_resp_bits_tagRdVec_5),
    .io_read_resp_bits_tagRdVec_6(dir_io_read_resp_bits_tagRdVec_6),
    .io_read_resp_bits_tagRdVec_7(dir_io_read_resp_bits_tagRdVec_7),
    .io_write_req_ready(dir_io_write_req_ready),
    .io_write_req_valid(dir_io_write_req_valid),
    .io_write_req_bits_addr(dir_io_write_req_bits_addr),
    .io_write_req_bits_way(dir_io_write_req_bits_way),
    .io_write_req_bits_meta(dir_io_write_req_bits_meta)
  );
  Arbiter mshrReqArb ( // @[DCache.scala 105:28]
    .io_in_0_ready(mshrReqArb_io_in_0_ready),
    .io_in_0_valid(mshrReqArb_io_in_0_valid),
    .io_in_0_bits_addr(mshrReqArb_io_in_0_bits_addr),
    .io_in_0_bits_dirInfo_hit(mshrReqArb_io_in_0_bits_dirInfo_hit),
    .io_in_0_bits_dirInfo_chosenWay(mshrReqArb_io_in_0_bits_dirInfo_chosenWay),
    .io_in_0_bits_dirInfo_isDirtyWay(mshrReqArb_io_in_0_bits_dirInfo_isDirtyWay),
    .io_in_0_bits_dirtyTag(mshrReqArb_io_in_0_bits_dirtyTag),
    .io_in_0_bits_data_0(mshrReqArb_io_in_0_bits_data_0),
    .io_in_0_bits_data_1(mshrReqArb_io_in_0_bits_data_1),
    .io_in_0_bits_data_2(mshrReqArb_io_in_0_bits_data_2),
    .io_in_0_bits_data_3(mshrReqArb_io_in_0_bits_data_3),
    .io_in_1_ready(mshrReqArb_io_in_1_ready),
    .io_in_1_valid(mshrReqArb_io_in_1_valid),
    .io_in_1_bits_addr(mshrReqArb_io_in_1_bits_addr),
    .io_in_1_bits_dirInfo_hit(mshrReqArb_io_in_1_bits_dirInfo_hit),
    .io_in_1_bits_dirInfo_chosenWay(mshrReqArb_io_in_1_bits_dirInfo_chosenWay),
    .io_in_1_bits_dirInfo_isDirtyWay(mshrReqArb_io_in_1_bits_dirInfo_isDirtyWay),
    .io_in_1_bits_dirtyTag(mshrReqArb_io_in_1_bits_dirtyTag),
    .io_in_1_bits_data_0(mshrReqArb_io_in_1_bits_data_0),
    .io_in_1_bits_data_1(mshrReqArb_io_in_1_bits_data_1),
    .io_in_1_bits_data_2(mshrReqArb_io_in_1_bits_data_2),
    .io_in_1_bits_data_3(mshrReqArb_io_in_1_bits_data_3),
    .io_in_1_bits_storeData(mshrReqArb_io_in_1_bits_storeData),
    .io_in_1_bits_storeMask(mshrReqArb_io_in_1_bits_storeMask),
    .io_out_ready(mshrReqArb_io_out_ready),
    .io_out_valid(mshrReqArb_io_out_valid),
    .io_out_bits_addr(mshrReqArb_io_out_bits_addr),
    .io_out_bits_dirInfo_hit(mshrReqArb_io_out_bits_dirInfo_hit),
    .io_out_bits_dirInfo_chosenWay(mshrReqArb_io_out_bits_dirInfo_chosenWay),
    .io_out_bits_dirInfo_isDirtyWay(mshrReqArb_io_out_bits_dirInfo_isDirtyWay),
    .io_out_bits_dirtyTag(mshrReqArb_io_out_bits_dirtyTag),
    .io_out_bits_data_0(mshrReqArb_io_out_bits_data_0),
    .io_out_bits_data_1(mshrReqArb_io_out_bits_data_1),
    .io_out_bits_data_2(mshrReqArb_io_out_bits_data_2),
    .io_out_bits_data_3(mshrReqArb_io_out_bits_data_3),
    .io_out_bits_isStore(mshrReqArb_io_out_bits_isStore),
    .io_out_bits_storeData(mshrReqArb_io_out_bits_storeData),
    .io_out_bits_storeMask(mshrReqArb_io_out_bits_storeMask)
  );
  Arbiter_1 tlbusReqArb ( // @[DCache.scala 110:29]
    .io_in_0_ready(tlbusReqArb_io_in_0_ready),
    .io_in_0_valid(tlbusReqArb_io_in_0_valid),
    .io_in_0_bits_address(tlbusReqArb_io_in_0_bits_address),
    .io_in_0_bits_data(tlbusReqArb_io_in_0_bits_data),
    .io_in_1_ready(tlbusReqArb_io_in_1_ready),
    .io_in_1_valid(tlbusReqArb_io_in_1_valid),
    .io_in_1_bits_address(tlbusReqArb_io_in_1_bits_address),
    .io_out_ready(tlbusReqArb_io_out_ready),
    .io_out_valid(tlbusReqArb_io_out_valid),
    .io_out_bits_opcode(tlbusReqArb_io_out_bits_opcode),
    .io_out_bits_address(tlbusReqArb_io_out_bits_address),
    .io_out_bits_data(tlbusReqArb_io_out_bits_data)
  );
  Arbiter_2 loadRespArb ( // @[DCache.scala 122:29]
    .io_in_0_valid(loadRespArb_io_in_0_valid),
    .io_in_0_bits_data(loadRespArb_io_in_0_bits_data),
    .io_in_1_ready(loadRespArb_io_in_1_ready),
    .io_in_1_valid(loadRespArb_io_in_1_valid),
    .io_in_1_bits_data(loadRespArb_io_in_1_bits_data),
    .io_out_valid(loadRespArb_io_out_valid),
    .io_out_bits_data(loadRespArb_io_out_bits_data)
  );
  Arbiter_3 storeRespArb ( // @[DCache.scala 127:30]
    .io_in_0_valid(storeRespArb_io_in_0_valid),
    .io_in_1_ready(storeRespArb_io_in_1_ready),
    .io_in_1_valid(storeRespArb_io_in_1_valid),
    .io_out_valid(storeRespArb_io_out_valid)
  );
  Arbiter_4 dbRdReqArb ( // @[DCache.scala 133:28]
    .io_in_0_valid(dbRdReqArb_io_in_0_valid),
    .io_in_0_bits_set(dbRdReqArb_io_in_0_bits_set),
    .io_in_1_ready(dbRdReqArb_io_in_1_ready),
    .io_in_1_valid(dbRdReqArb_io_in_1_valid),
    .io_in_1_bits_set(dbRdReqArb_io_in_1_bits_set),
    .io_out_valid(dbRdReqArb_io_out_valid),
    .io_out_bits_set(dbRdReqArb_io_out_bits_set)
  );
  Arbiter_5 dirRdReqArb ( // @[DCache.scala 138:29]
    .io_in_0_valid(dirRdReqArb_io_in_0_valid),
    .io_in_0_bits_addr(dirRdReqArb_io_in_0_bits_addr),
    .io_in_1_ready(dirRdReqArb_io_in_1_ready),
    .io_in_1_valid(dirRdReqArb_io_in_1_valid),
    .io_in_1_bits_addr(dirRdReqArb_io_in_1_bits_addr),
    .io_out_valid(dirRdReqArb_io_out_valid),
    .io_out_bits_addr(dirRdReqArb_io_out_bits_addr)
  );
  Arbiter_6 dataBankWrArb ( // @[DCache.scala 144:31]
    .io_in_0_valid(dataBankWrArb_io_in_0_valid),
    .io_in_0_bits_set(dataBankWrArb_io_in_0_bits_set),
    .io_in_0_bits_data_0(dataBankWrArb_io_in_0_bits_data_0),
    .io_in_0_bits_data_1(dataBankWrArb_io_in_0_bits_data_1),
    .io_in_0_bits_data_2(dataBankWrArb_io_in_0_bits_data_2),
    .io_in_0_bits_data_3(dataBankWrArb_io_in_0_bits_data_3),
    .io_in_0_bits_blockMask(dataBankWrArb_io_in_0_bits_blockMask),
    .io_in_0_bits_way(dataBankWrArb_io_in_0_bits_way),
    .io_in_1_ready(dataBankWrArb_io_in_1_ready),
    .io_in_1_valid(dataBankWrArb_io_in_1_valid),
    .io_in_1_bits_set(dataBankWrArb_io_in_1_bits_set),
    .io_in_1_bits_data_0(dataBankWrArb_io_in_1_bits_data_0),
    .io_in_1_bits_data_1(dataBankWrArb_io_in_1_bits_data_1),
    .io_in_1_bits_data_2(dataBankWrArb_io_in_1_bits_data_2),
    .io_in_1_bits_data_3(dataBankWrArb_io_in_1_bits_data_3),
    .io_in_1_bits_way(dataBankWrArb_io_in_1_bits_way),
    .io_in_2_ready(dataBankWrArb_io_in_2_ready),
    .io_in_2_valid(dataBankWrArb_io_in_2_valid),
    .io_in_2_bits_set(dataBankWrArb_io_in_2_bits_set),
    .io_in_2_bits_data_0(dataBankWrArb_io_in_2_bits_data_0),
    .io_in_2_bits_data_1(dataBankWrArb_io_in_2_bits_data_1),
    .io_in_2_bits_data_2(dataBankWrArb_io_in_2_bits_data_2),
    .io_in_2_bits_data_3(dataBankWrArb_io_in_2_bits_data_3),
    .io_in_2_bits_blockMask(dataBankWrArb_io_in_2_bits_blockMask),
    .io_in_2_bits_way(dataBankWrArb_io_in_2_bits_way),
    .io_out_valid(dataBankWrArb_io_out_valid),
    .io_out_bits_set(dataBankWrArb_io_out_bits_set),
    .io_out_bits_data_0(dataBankWrArb_io_out_bits_data_0),
    .io_out_bits_data_1(dataBankWrArb_io_out_bits_data_1),
    .io_out_bits_data_2(dataBankWrArb_io_out_bits_data_2),
    .io_out_bits_data_3(dataBankWrArb_io_out_bits_data_3),
    .io_out_bits_blockMask(dataBankWrArb_io_out_bits_blockMask),
    .io_out_bits_way(dataBankWrArb_io_out_bits_way)
  );
  Arbiter_7 dirWrArb ( // @[DCache.scala 150:26]
    .io_in_0_valid(dirWrArb_io_in_0_valid),
    .io_in_0_bits_addr(dirWrArb_io_in_0_bits_addr),
    .io_in_0_bits_way(dirWrArb_io_in_0_bits_way),
    .io_in_1_ready(dirWrArb_io_in_1_ready),
    .io_in_1_valid(dirWrArb_io_in_1_valid),
    .io_in_1_bits_addr(dirWrArb_io_in_1_bits_addr),
    .io_in_1_bits_way(dirWrArb_io_in_1_bits_way),
    .io_in_2_ready(dirWrArb_io_in_2_ready),
    .io_in_2_valid(dirWrArb_io_in_2_valid),
    .io_in_2_bits_addr(dirWrArb_io_in_2_bits_addr),
    .io_in_2_bits_way(dirWrArb_io_in_2_bits_way),
    .io_out_valid(dirWrArb_io_out_valid),
    .io_out_bits_addr(dirWrArb_io_out_bits_addr),
    .io_out_bits_way(dirWrArb_io_out_bits_way),
    .io_out_bits_meta(dirWrArb_io_out_bits_meta)
  );
  assign io_read_req_ready = loadPipe_io_load_req_ready; // @[DCache.scala 97:26]
  assign io_read_resp_valid = loadRespArb_io_out_valid; // @[DCache.scala 125:18]
  assign io_read_resp_bits_data = loadRespArb_io_out_bits_data; // @[DCache.scala 125:18]
  assign io_write_req_ready = storePipe_io_store_req_ready; // @[DCache.scala 98:28]
  assign io_write_resp_valid = storeRespArb_io_out_valid; // @[DCache.scala 130:19]
  assign io_tlbus_req_valid = tlbusReqArb_io_out_valid; // @[DCache.scala 113:18]
  assign io_tlbus_req_bits_opcode = tlbusReqArb_io_out_bits_opcode; // @[DCache.scala 113:18]
  assign io_tlbus_req_bits_address = tlbusReqArb_io_out_bits_address; // @[DCache.scala 113:18]
  assign io_tlbus_req_bits_data = tlbusReqArb_io_out_bits_data; // @[DCache.scala 113:18]
  assign io_tlbus_resp_ready = 1'h1; // @[DCache.scala 119:51]
  assign loadPipe_clock = clock;
  assign loadPipe_reset = reset;
  assign loadPipe_io_load_req_valid = io_read_req_valid; // @[DCache.scala 97:26]
  assign loadPipe_io_load_req_bits_addr = io_read_req_bits_addr; // @[DCache.scala 97:26]
  assign loadPipe_io_dir_req_ready = dirRdReqArb_io_in_1_ready; // @[DCache.scala 140:26]
  assign loadPipe_io_dir_resp_bits_hit = dir_io_read_resp_bits_hit; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_chosenWay = dir_io_read_resp_bits_chosenWay; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_isDirtyWay = dir_io_read_resp_bits_isDirtyWay; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_0 = dir_io_read_resp_bits_tagRdVec_0; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_1 = dir_io_read_resp_bits_tagRdVec_1; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_2 = dir_io_read_resp_bits_tagRdVec_2; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_3 = dir_io_read_resp_bits_tagRdVec_3; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_4 = dir_io_read_resp_bits_tagRdVec_4; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_5 = dir_io_read_resp_bits_tagRdVec_5; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_6 = dir_io_read_resp_bits_tagRdVec_6; // @[DCache.scala 90:31]
  assign loadPipe_io_dir_resp_bits_tagRdVec_7 = dir_io_read_resp_bits_tagRdVec_7; // @[DCache.scala 90:31]
  assign loadPipe_io_dataBank_req_ready = dbRdReqArb_io_in_1_ready; // @[DCache.scala 135:25]
  assign loadPipe_io_dataBank_resp_0_0 = db_io_read_resp_0_0; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_0_1 = db_io_read_resp_0_1; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_0_2 = db_io_read_resp_0_2; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_0_3 = db_io_read_resp_0_3; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_1_0 = db_io_read_resp_1_0; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_1_1 = db_io_read_resp_1_1; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_1_2 = db_io_read_resp_1_2; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_1_3 = db_io_read_resp_1_3; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_2_0 = db_io_read_resp_2_0; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_2_1 = db_io_read_resp_2_1; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_2_2 = db_io_read_resp_2_2; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_2_3 = db_io_read_resp_2_3; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_3_0 = db_io_read_resp_3_0; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_3_1 = db_io_read_resp_3_1; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_3_2 = db_io_read_resp_3_2; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_3_3 = db_io_read_resp_3_3; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_4_0 = db_io_read_resp_4_0; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_4_1 = db_io_read_resp_4_1; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_4_2 = db_io_read_resp_4_2; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_4_3 = db_io_read_resp_4_3; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_5_0 = db_io_read_resp_5_0; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_5_1 = db_io_read_resp_5_1; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_5_2 = db_io_read_resp_5_2; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_5_3 = db_io_read_resp_5_3; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_6_0 = db_io_read_resp_6_0; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_6_1 = db_io_read_resp_6_1; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_6_2 = db_io_read_resp_6_2; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_6_3 = db_io_read_resp_6_3; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_7_0 = db_io_read_resp_7_0; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_7_1 = db_io_read_resp_7_1; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_7_2 = db_io_read_resp_7_2; // @[DCache.scala 94:31]
  assign loadPipe_io_dataBank_resp_7_3 = db_io_read_resp_7_3; // @[DCache.scala 94:31]
  assign loadPipe_io_mshr_ready = mshrReqArb_io_in_0_ready; // @[DCache.scala 106:25]
  assign storePipe_clock = clock;
  assign storePipe_reset = reset;
  assign storePipe_io_store_req_valid = io_write_req_valid; // @[DCache.scala 98:28]
  assign storePipe_io_store_req_bits_addr = io_write_req_bits_addr; // @[DCache.scala 98:28]
  assign storePipe_io_store_req_bits_data = io_write_req_bits_data; // @[DCache.scala 98:28]
  assign storePipe_io_store_req_bits_mask = io_write_req_bits_mask; // @[DCache.scala 98:28]
  assign storePipe_io_dir_read_resp_bits_hit = dir_io_read_resp_bits_hit; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_chosenWay = dir_io_read_resp_bits_chosenWay; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_isDirtyWay = dir_io_read_resp_bits_isDirtyWay; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_0 = dir_io_read_resp_bits_tagRdVec_0; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_1 = dir_io_read_resp_bits_tagRdVec_1; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_2 = dir_io_read_resp_bits_tagRdVec_2; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_3 = dir_io_read_resp_bits_tagRdVec_3; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_4 = dir_io_read_resp_bits_tagRdVec_4; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_5 = dir_io_read_resp_bits_tagRdVec_5; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_6 = dir_io_read_resp_bits_tagRdVec_6; // @[DCache.scala 92:37]
  assign storePipe_io_dir_read_resp_bits_tagRdVec_7 = dir_io_read_resp_bits_tagRdVec_7; // @[DCache.scala 92:37]
  assign storePipe_io_dataBank_read_resp_0_0 = db_io_read_resp_0_0; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_0_1 = db_io_read_resp_0_1; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_0_2 = db_io_read_resp_0_2; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_0_3 = db_io_read_resp_0_3; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_1_0 = db_io_read_resp_1_0; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_1_1 = db_io_read_resp_1_1; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_1_2 = db_io_read_resp_1_2; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_1_3 = db_io_read_resp_1_3; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_2_0 = db_io_read_resp_2_0; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_2_1 = db_io_read_resp_2_1; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_2_2 = db_io_read_resp_2_2; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_2_3 = db_io_read_resp_2_3; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_3_0 = db_io_read_resp_3_0; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_3_1 = db_io_read_resp_3_1; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_3_2 = db_io_read_resp_3_2; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_3_3 = db_io_read_resp_3_3; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_4_0 = db_io_read_resp_4_0; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_4_1 = db_io_read_resp_4_1; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_4_2 = db_io_read_resp_4_2; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_4_3 = db_io_read_resp_4_3; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_5_0 = db_io_read_resp_5_0; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_5_1 = db_io_read_resp_5_1; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_5_2 = db_io_read_resp_5_2; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_5_3 = db_io_read_resp_5_3; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_6_0 = db_io_read_resp_6_0; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_6_1 = db_io_read_resp_6_1; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_6_2 = db_io_read_resp_6_2; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_6_3 = db_io_read_resp_6_3; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_7_0 = db_io_read_resp_7_0; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_7_1 = db_io_read_resp_7_1; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_7_2 = db_io_read_resp_7_2; // @[DCache.scala 95:37]
  assign storePipe_io_dataBank_read_resp_7_3 = db_io_read_resp_7_3; // @[DCache.scala 95:37]
  assign storePipe_io_mshr_ready = mshrReqArb_io_in_1_ready; // @[DCache.scala 107:25]
  assign mshr_clock = clock;
  assign mshr_reset = reset;
  assign mshr_io_req_valid = mshrReqArb_io_out_valid; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_addr = mshrReqArb_io_out_bits_addr; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_dirInfo_hit = mshrReqArb_io_out_bits_dirInfo_hit; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_dirInfo_chosenWay = mshrReqArb_io_out_bits_dirInfo_chosenWay; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_dirInfo_isDirtyWay = mshrReqArb_io_out_bits_dirInfo_isDirtyWay; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_dirtyTag = mshrReqArb_io_out_bits_dirtyTag; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_data_0 = mshrReqArb_io_out_bits_data_0; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_data_1 = mshrReqArb_io_out_bits_data_1; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_data_2 = mshrReqArb_io_out_bits_data_2; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_data_3 = mshrReqArb_io_out_bits_data_3; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_isStore = mshrReqArb_io_out_bits_isStore; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_storeData = mshrReqArb_io_out_bits_storeData; // @[DCache.scala 108:17]
  assign mshr_io_req_bits_storeMask = mshrReqArb_io_out_bits_storeMask; // @[DCache.scala 108:17]
  assign mshr_io_resp_load_ready = loadRespArb_io_in_1_ready; // @[DCache.scala 124:26]
  assign mshr_io_resp_store_ready = storeRespArb_io_in_1_ready; // @[DCache.scala 129:27]
  assign mshr_io_tasks_refill_resp_valid = refillPipe_io_resp_valid; // @[DCache.scala 101:31]
  assign mshr_io_tasks_refill_resp_bits_data = refillPipe_io_resp_bits_data; // @[DCache.scala 101:31]
  assign mshr_io_tasks_writeback_resp_valid = wb_io_resp_valid; // @[DCache.scala 103:34]
  assign mshr_io_dirWrite_req_ready = dirWrArb_io_in_2_ready; // @[DCache.scala 153:23]
  assign mshr_io_dataWrite_req_ready = dataBankWrArb_io_in_2_ready; // @[DCache.scala 147:28]
  assign refillPipe_clock = clock;
  assign refillPipe_reset = reset;
  assign refillPipe_io_req_valid = mshr_io_tasks_refill_req_valid; // @[DCache.scala 100:30]
  assign refillPipe_io_req_bits_addr = mshr_io_tasks_refill_req_bits_addr; // @[DCache.scala 100:30]
  assign refillPipe_io_req_bits_chosenWay = mshr_io_tasks_refill_req_bits_chosenWay; // @[DCache.scala 100:30]
  assign refillPipe_io_tlbus_req_ready = tlbusReqArb_io_in_1_ready; // @[DCache.scala 112:26]
  assign refillPipe_io_tlbus_resp_valid = io_tlbus_resp_valid; // @[DCache.scala 117:36]
  assign refillPipe_io_tlbus_resp_bits_opcode = io_tlbus_resp_bits_opcode; // @[DCache.scala 118:35]
  assign refillPipe_io_tlbus_resp_bits_data = io_tlbus_resp_bits_data; // @[DCache.scala 118:35]
  assign refillPipe_io_dirWrite_req_ready = dirWrArb_io_in_1_ready; // @[DCache.scala 152:23]
  assign refillPipe_io_dataWrite_req_ready = dataBankWrArb_io_in_1_ready; // @[DCache.scala 146:28]
  assign wb_clock = clock;
  assign wb_reset = reset;
  assign wb_io_req_valid = mshr_io_tasks_writeback_req_valid; // @[DCache.scala 102:33]
  assign wb_io_req_bits_addr = mshr_io_tasks_writeback_req_bits_addr; // @[DCache.scala 102:33]
  assign wb_io_req_bits_dirtyTag = mshr_io_tasks_writeback_req_bits_dirtyTag; // @[DCache.scala 102:33]
  assign wb_io_req_bits_data_0 = mshr_io_tasks_writeback_req_bits_data_0; // @[DCache.scala 102:33]
  assign wb_io_req_bits_data_1 = mshr_io_tasks_writeback_req_bits_data_1; // @[DCache.scala 102:33]
  assign wb_io_req_bits_data_2 = mshr_io_tasks_writeback_req_bits_data_2; // @[DCache.scala 102:33]
  assign wb_io_req_bits_data_3 = mshr_io_tasks_writeback_req_bits_data_3; // @[DCache.scala 102:33]
  assign wb_io_tlbus_req_ready = tlbusReqArb_io_in_0_ready; // @[DCache.scala 111:26]
  assign wb_io_tlbus_resp_valid = io_tlbus_resp_valid; // @[DCache.scala 115:28]
  assign db_clock = clock;
  assign db_reset = reset;
  assign db_io_read_req_valid = dbRdReqArb_io_out_valid; // @[DCache.scala 136:20]
  assign db_io_read_req_bits_set = dbRdReqArb_io_out_bits_set; // @[DCache.scala 136:20]
  assign db_io_write_req_valid = dataBankWrArb_io_out_valid; // @[DCache.scala 148:21]
  assign db_io_write_req_bits_set = dataBankWrArb_io_out_bits_set; // @[DCache.scala 148:21]
  assign db_io_write_req_bits_data_0 = dataBankWrArb_io_out_bits_data_0; // @[DCache.scala 148:21]
  assign db_io_write_req_bits_data_1 = dataBankWrArb_io_out_bits_data_1; // @[DCache.scala 148:21]
  assign db_io_write_req_bits_data_2 = dataBankWrArb_io_out_bits_data_2; // @[DCache.scala 148:21]
  assign db_io_write_req_bits_data_3 = dataBankWrArb_io_out_bits_data_3; // @[DCache.scala 148:21]
  assign db_io_write_req_bits_blockMask = dataBankWrArb_io_out_bits_blockMask; // @[DCache.scala 148:21]
  assign db_io_write_req_bits_way = dataBankWrArb_io_out_bits_way; // @[DCache.scala 148:21]
  assign dir_clock = clock;
  assign dir_reset = reset;
  assign dir_io_read_req_valid = dirRdReqArb_io_out_valid; // @[DCache.scala 141:21]
  assign dir_io_read_req_bits_addr = dirRdReqArb_io_out_bits_addr; // @[DCache.scala 141:21]
  assign dir_io_write_req_valid = dirWrArb_io_out_valid; // @[DCache.scala 154:22]
  assign dir_io_write_req_bits_addr = dirWrArb_io_out_bits_addr; // @[DCache.scala 154:22]
  assign dir_io_write_req_bits_way = dirWrArb_io_out_bits_way; // @[DCache.scala 154:22]
  assign dir_io_write_req_bits_meta = dirWrArb_io_out_bits_meta; // @[DCache.scala 154:22]
  assign mshrReqArb_io_in_0_valid = loadPipe_io_mshr_valid; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_0_bits_addr = loadPipe_io_mshr_bits_addr; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_0_bits_dirInfo_hit = loadPipe_io_mshr_bits_dirInfo_hit; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_0_bits_dirInfo_chosenWay = loadPipe_io_mshr_bits_dirInfo_chosenWay; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_0_bits_dirInfo_isDirtyWay = loadPipe_io_mshr_bits_dirInfo_isDirtyWay; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_0_bits_dirtyTag = loadPipe_io_mshr_bits_dirtyTag; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_0_bits_data_0 = loadPipe_io_mshr_bits_data_0; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_0_bits_data_1 = loadPipe_io_mshr_bits_data_1; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_0_bits_data_2 = loadPipe_io_mshr_bits_data_2; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_0_bits_data_3 = loadPipe_io_mshr_bits_data_3; // @[DCache.scala 106:25]
  assign mshrReqArb_io_in_1_valid = storePipe_io_mshr_valid; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_addr = storePipe_io_mshr_bits_addr; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_dirInfo_hit = storePipe_io_mshr_bits_dirInfo_hit; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_dirInfo_chosenWay = storePipe_io_mshr_bits_dirInfo_chosenWay; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_dirInfo_isDirtyWay = storePipe_io_mshr_bits_dirInfo_isDirtyWay; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_dirtyTag = storePipe_io_mshr_bits_dirtyTag; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_data_0 = storePipe_io_mshr_bits_data_0; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_data_1 = storePipe_io_mshr_bits_data_1; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_data_2 = storePipe_io_mshr_bits_data_2; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_data_3 = storePipe_io_mshr_bits_data_3; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_storeData = storePipe_io_mshr_bits_storeData; // @[DCache.scala 107:25]
  assign mshrReqArb_io_in_1_bits_storeMask = storePipe_io_mshr_bits_storeMask; // @[DCache.scala 107:25]
  assign mshrReqArb_io_out_ready = mshr_io_req_ready; // @[DCache.scala 108:17]
  assign tlbusReqArb_io_in_0_valid = wb_io_tlbus_req_valid; // @[DCache.scala 111:26]
  assign tlbusReqArb_io_in_0_bits_address = wb_io_tlbus_req_bits_address; // @[DCache.scala 111:26]
  assign tlbusReqArb_io_in_0_bits_data = wb_io_tlbus_req_bits_data; // @[DCache.scala 111:26]
  assign tlbusReqArb_io_in_1_valid = refillPipe_io_tlbus_req_valid; // @[DCache.scala 112:26]
  assign tlbusReqArb_io_in_1_bits_address = refillPipe_io_tlbus_req_bits_address; // @[DCache.scala 112:26]
  assign tlbusReqArb_io_out_ready = io_tlbus_req_ready; // @[DCache.scala 113:18]
  assign loadRespArb_io_in_0_valid = loadPipe_io_load_resp_valid; // @[DCache.scala 123:26]
  assign loadRespArb_io_in_0_bits_data = loadPipe_io_load_resp_bits_data; // @[DCache.scala 123:26]
  assign loadRespArb_io_in_1_valid = mshr_io_resp_load_valid; // @[DCache.scala 124:26]
  assign loadRespArb_io_in_1_bits_data = mshr_io_resp_load_bits_data; // @[DCache.scala 124:26]
  assign storeRespArb_io_in_0_valid = storePipe_io_store_resp_valid; // @[DCache.scala 128:27]
  assign storeRespArb_io_in_1_valid = mshr_io_resp_store_valid; // @[DCache.scala 129:27]
  assign dbRdReqArb_io_in_0_valid = storePipe_io_dataBank_read_req_valid; // @[DCache.scala 134:25]
  assign dbRdReqArb_io_in_0_bits_set = storePipe_io_dataBank_read_req_bits_set; // @[DCache.scala 134:25]
  assign dbRdReqArb_io_in_1_valid = loadPipe_io_dataBank_req_valid; // @[DCache.scala 135:25]
  assign dbRdReqArb_io_in_1_bits_set = loadPipe_io_dataBank_req_bits_set; // @[DCache.scala 135:25]
  assign dirRdReqArb_io_in_0_valid = storePipe_io_dir_read_req_valid; // @[DCache.scala 139:26]
  assign dirRdReqArb_io_in_0_bits_addr = storePipe_io_dir_read_req_bits_addr; // @[DCache.scala 139:26]
  assign dirRdReqArb_io_in_1_valid = loadPipe_io_dir_req_valid; // @[DCache.scala 140:26]
  assign dirRdReqArb_io_in_1_bits_addr = loadPipe_io_dir_req_bits_addr; // @[DCache.scala 140:26]
  assign dataBankWrArb_io_in_0_valid = storePipe_io_dataBank_write_req_valid; // @[DCache.scala 145:28]
  assign dataBankWrArb_io_in_0_bits_set = storePipe_io_dataBank_write_req_bits_set; // @[DCache.scala 145:28]
  assign dataBankWrArb_io_in_0_bits_data_0 = storePipe_io_dataBank_write_req_bits_data_0; // @[DCache.scala 145:28]
  assign dataBankWrArb_io_in_0_bits_data_1 = storePipe_io_dataBank_write_req_bits_data_1; // @[DCache.scala 145:28]
  assign dataBankWrArb_io_in_0_bits_data_2 = storePipe_io_dataBank_write_req_bits_data_2; // @[DCache.scala 145:28]
  assign dataBankWrArb_io_in_0_bits_data_3 = storePipe_io_dataBank_write_req_bits_data_3; // @[DCache.scala 145:28]
  assign dataBankWrArb_io_in_0_bits_blockMask = storePipe_io_dataBank_write_req_bits_blockMask; // @[DCache.scala 145:28]
  assign dataBankWrArb_io_in_0_bits_way = storePipe_io_dataBank_write_req_bits_way; // @[DCache.scala 145:28]
  assign dataBankWrArb_io_in_1_valid = refillPipe_io_dataWrite_req_valid; // @[DCache.scala 146:28]
  assign dataBankWrArb_io_in_1_bits_set = refillPipe_io_dataWrite_req_bits_set; // @[DCache.scala 146:28]
  assign dataBankWrArb_io_in_1_bits_data_0 = refillPipe_io_dataWrite_req_bits_data_0; // @[DCache.scala 146:28]
  assign dataBankWrArb_io_in_1_bits_data_1 = refillPipe_io_dataWrite_req_bits_data_1; // @[DCache.scala 146:28]
  assign dataBankWrArb_io_in_1_bits_data_2 = refillPipe_io_dataWrite_req_bits_data_2; // @[DCache.scala 146:28]
  assign dataBankWrArb_io_in_1_bits_data_3 = refillPipe_io_dataWrite_req_bits_data_3; // @[DCache.scala 146:28]
  assign dataBankWrArb_io_in_1_bits_way = refillPipe_io_dataWrite_req_bits_way; // @[DCache.scala 146:28]
  assign dataBankWrArb_io_in_2_valid = mshr_io_dataWrite_req_valid; // @[DCache.scala 147:28]
  assign dataBankWrArb_io_in_2_bits_set = mshr_io_dataWrite_req_bits_set; // @[DCache.scala 147:28]
  assign dataBankWrArb_io_in_2_bits_data_0 = mshr_io_dataWrite_req_bits_data_0; // @[DCache.scala 147:28]
  assign dataBankWrArb_io_in_2_bits_data_1 = mshr_io_dataWrite_req_bits_data_1; // @[DCache.scala 147:28]
  assign dataBankWrArb_io_in_2_bits_data_2 = mshr_io_dataWrite_req_bits_data_2; // @[DCache.scala 147:28]
  assign dataBankWrArb_io_in_2_bits_data_3 = mshr_io_dataWrite_req_bits_data_3; // @[DCache.scala 147:28]
  assign dataBankWrArb_io_in_2_bits_blockMask = mshr_io_dataWrite_req_bits_blockMask; // @[DCache.scala 147:28]
  assign dataBankWrArb_io_in_2_bits_way = mshr_io_dataWrite_req_bits_way; // @[DCache.scala 147:28]
  assign dirWrArb_io_in_0_valid = storePipe_io_dir_write_req_valid; // @[DCache.scala 151:23]
  assign dirWrArb_io_in_0_bits_addr = storePipe_io_dir_write_req_bits_addr; // @[DCache.scala 151:23]
  assign dirWrArb_io_in_0_bits_way = storePipe_io_dir_write_req_bits_way; // @[DCache.scala 151:23]
  assign dirWrArb_io_in_1_valid = refillPipe_io_dirWrite_req_valid; // @[DCache.scala 152:23]
  assign dirWrArb_io_in_1_bits_addr = refillPipe_io_dirWrite_req_bits_addr; // @[DCache.scala 152:23]
  assign dirWrArb_io_in_1_bits_way = refillPipe_io_dirWrite_req_bits_way; // @[DCache.scala 152:23]
  assign dirWrArb_io_in_2_valid = mshr_io_dirWrite_req_valid; // @[DCache.scala 153:23]
  assign dirWrArb_io_in_2_bits_addr = mshr_io_dirWrite_req_bits_addr; // @[DCache.scala 153:23]
  assign dirWrArb_io_in_2_bits_way = mshr_io_dirWrite_req_bits_way; // @[DCache.scala 153:23]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 162:24]
      c <= 64'h0; // @[util.scala 162:24]
    end else begin
      c <= _c_T_1; // @[util.scala 163:11]
    end
    if (reset) begin // @[util.scala 162:24]
      c_1 <= 64'h0; // @[util.scala 162:24]
    end else begin
      c_1 <= _c_T_3; // @[util.scala 163:11]
    end
    if (reset) begin // @[util.scala 162:24]
      c_2 <= 64'h0; // @[util.scala 162:24]
    end else begin
      c_2 <= _c_T_5; // @[util.scala 163:11]
    end
    if (reset) begin // @[util.scala 162:24]
      c_3 <= 64'h0; // @[util.scala 162:24]
    end else begin
      c_3 <= _c_T_7; // @[util.scala 163:11]
    end
    if (reset) begin // @[util.scala 162:24]
      c_4 <= 64'h0; // @[util.scala 162:24]
    end else begin
      c_4 <= _c_T_9; // @[util.scala 163:11]
    end
    if (reset) begin // @[util.scala 162:24]
      c_5 <= 64'h0; // @[util.scala 162:24]
    end else begin
      c_5 <= _c_T_11; // @[util.scala 163:11]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [DCache] read req ==> addr: 0x%x\n",c,io_read_req_bits_addr); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_read_resp_valid & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [DCache] read resp <== data: 0x%x\n",c_1,io_read_resp_bits_data); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [DCache] write req ==> addr: 0x%x  data: 0x%x\n",c_2,
            io_write_req_bits_addr,io_write_req_bits_data); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_write_resp_valid & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [DCache] write resp <== \n",c_3); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14 & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [DCache] dirty write back ==> data: 0x%x  addr: 0x%x\n",c_4,
            io_tlbus_req_bits_data,io_tlbus_req_bits_address); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_19 & ~reset) begin
          $fwrite(32'h80000002,"[SimLog ][time=%d] [DCache] refill resp <== data: 0x%x ",c_5,io_tlbus_resp_bits_data); // @[util.scala 16:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  c_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  c_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  c_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  c_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c_5 = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Mem(
  input          clock,
  input          reset,
  output         io_in_ready,
  input  [1:0]   io_in_bits_resultSrc,
  input  [4:0]   io_in_bits_lsuOp,
  input          io_in_bits_regWrEn,
  input  [31:0]  io_in_bits_aluOut,
  input  [31:0]  io_in_bits_data2,
  input  [31:0]  io_in_bits_pcNext4,
  input  [2:0]   io_in_bits_csrOp,
  input          io_in_bits_csrWrEn,
  input          io_in_bits_csrValid,
  input  [31:0]  io_in_bits_csrRdData,
  input  [31:0]  io_in_bits_csrWrData,
  input  [31:0]  io_in_bits_csrAddr,
  input  [3:0]   io_in_bits_excType,
  input          io_in_bits_instState_commit,
  input  [31:0]  io_in_bits_instState_pc,
  input  [31:0]  io_in_bits_instState_inst,
  input          io_out_ready,
  output         io_out_valid,
  output [1:0]   io_out_bits_resultSrc,
  output         io_out_bits_regWrEn,
  output [31:0]  io_out_bits_aluOut,
  output [31:0]  io_out_bits_pcNext4,
  output [2:0]   io_out_bits_csrOp,
  output         io_out_bits_csrWrEn,
  output [31:0]  io_out_bits_csrRdData,
  output [31:0]  io_out_bits_csrWrData,
  output [11:0]  io_out_bits_csrAddr,
  output         io_out_bits_instState_commit,
  output [31:0]  io_out_bits_instState_pc,
  output [31:0]  io_out_bits_instState_inst,
  output [31:0]  io_lsuData,
  output         io_lsuOK,
  input          io_tlbus_req_ready,
  output         io_tlbus_req_valid,
  output [2:0]   io_tlbus_req_bits_opcode,
  output [31:0]  io_tlbus_req_bits_address,
  output [127:0] io_tlbus_req_bits_data,
  input          io_tlbus_resp_valid,
  input  [2:0]   io_tlbus_resp_bits_opcode,
  input  [127:0] io_tlbus_resp_bits_data,
  output [4:0]   io_hazard_rd,
  output [31:0]  io_hazard_rdVal,
  output         io_hazard_regWrEn,
  input          io_ctrl_flush,
  output         io_excp_valid,
  output         io_excp_bits_isMret,
  output         io_excp_bits_isSret,
  output [30:0]  io_excp_bits_excCause,
  output [31:0]  io_excp_bits_excPc,
  input          io_csrBusy,
  input  [1:0]   io_csrMode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  lsu_clock; // @[4_Mem.scala 146:21]
  wire  lsu_reset; // @[4_Mem.scala 146:21]
  wire  lsu_io_req_ready; // @[4_Mem.scala 146:21]
  wire  lsu_io_req_valid; // @[4_Mem.scala 146:21]
  wire [31:0] lsu_io_req_bits_addr; // @[4_Mem.scala 146:21]
  wire [31:0] lsu_io_req_bits_wdata; // @[4_Mem.scala 146:21]
  wire [4:0] lsu_io_req_bits_lsuOp; // @[4_Mem.scala 146:21]
  wire  lsu_io_resp_valid; // @[4_Mem.scala 146:21]
  wire [31:0] lsu_io_resp_bits_rdata; // @[4_Mem.scala 146:21]
  wire  lsu_io_cache_read_req_ready; // @[4_Mem.scala 146:21]
  wire  lsu_io_cache_read_req_valid; // @[4_Mem.scala 146:21]
  wire [31:0] lsu_io_cache_read_req_bits_addr; // @[4_Mem.scala 146:21]
  wire  lsu_io_cache_read_resp_ready; // @[4_Mem.scala 146:21]
  wire  lsu_io_cache_read_resp_valid; // @[4_Mem.scala 146:21]
  wire [31:0] lsu_io_cache_read_resp_bits_data; // @[4_Mem.scala 146:21]
  wire  lsu_io_cache_write_req_ready; // @[4_Mem.scala 146:21]
  wire  lsu_io_cache_write_req_valid; // @[4_Mem.scala 146:21]
  wire [31:0] lsu_io_cache_write_req_bits_addr; // @[4_Mem.scala 146:21]
  wire [31:0] lsu_io_cache_write_req_bits_data; // @[4_Mem.scala 146:21]
  wire [3:0] lsu_io_cache_write_req_bits_mask; // @[4_Mem.scala 146:21]
  wire  lsu_io_cache_write_resp_ready; // @[4_Mem.scala 146:21]
  wire  lsu_io_cache_write_resp_valid; // @[4_Mem.scala 146:21]
  wire  dcache_clock; // @[4_Mem.scala 165:24]
  wire  dcache_reset; // @[4_Mem.scala 165:24]
  wire  dcache_io_read_req_ready; // @[4_Mem.scala 165:24]
  wire  dcache_io_read_req_valid; // @[4_Mem.scala 165:24]
  wire [31:0] dcache_io_read_req_bits_addr; // @[4_Mem.scala 165:24]
  wire  dcache_io_read_resp_valid; // @[4_Mem.scala 165:24]
  wire [31:0] dcache_io_read_resp_bits_data; // @[4_Mem.scala 165:24]
  wire  dcache_io_write_req_ready; // @[4_Mem.scala 165:24]
  wire  dcache_io_write_req_valid; // @[4_Mem.scala 165:24]
  wire [31:0] dcache_io_write_req_bits_addr; // @[4_Mem.scala 165:24]
  wire [31:0] dcache_io_write_req_bits_data; // @[4_Mem.scala 165:24]
  wire [3:0] dcache_io_write_req_bits_mask; // @[4_Mem.scala 165:24]
  wire  dcache_io_write_resp_valid; // @[4_Mem.scala 165:24]
  wire  dcache_io_tlbus_req_ready; // @[4_Mem.scala 165:24]
  wire  dcache_io_tlbus_req_valid; // @[4_Mem.scala 165:24]
  wire [2:0] dcache_io_tlbus_req_bits_opcode; // @[4_Mem.scala 165:24]
  wire [31:0] dcache_io_tlbus_req_bits_address; // @[4_Mem.scala 165:24]
  wire [127:0] dcache_io_tlbus_req_bits_data; // @[4_Mem.scala 165:24]
  wire  dcache_io_tlbus_resp_ready; // @[4_Mem.scala 165:24]
  wire  dcache_io_tlbus_resp_valid; // @[4_Mem.scala 165:24]
  wire [2:0] dcache_io_tlbus_resp_bits_opcode; // @[4_Mem.scala 165:24]
  wire [127:0] dcache_io_tlbus_resp_bits_data; // @[4_Mem.scala 165:24]
  wire  lsuReady = lsu_io_req_ready; // @[4_Mem.scala 148:14 60:28]
  reg [4:0] stageReg_lsuOp; // @[4_Mem.scala 70:27]
  wire  validLsuOp = ~(stageReg_lsuOp == 5'h0 | stageReg_lsuOp == 5'h14); // @[4_Mem.scala 149:19]
  wire  stall = ~lsuReady | validLsuOp & ~io_lsuOK; // @[4_Mem.scala 64:44]
  wire  _io_in_ready_T = ~stall; // @[4_Mem.scala 68:20]
  wire  _io_in_ready_T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  reg [1:0] stageReg_resultSrc; // @[4_Mem.scala 70:27]
  reg  stageReg_regWrEn; // @[4_Mem.scala 70:27]
  reg [31:0] stageReg_aluOut; // @[4_Mem.scala 70:27]
  reg [31:0] stageReg_data2; // @[4_Mem.scala 70:27]
  reg [31:0] stageReg_pcNext4; // @[4_Mem.scala 70:27]
  reg [2:0] stageReg_csrOp; // @[4_Mem.scala 70:27]
  reg  stageReg_csrWrEn; // @[4_Mem.scala 70:27]
  reg  stageReg_csrValid; // @[4_Mem.scala 70:27]
  reg [31:0] stageReg_csrRdData; // @[4_Mem.scala 70:27]
  reg [31:0] stageReg_csrWrData; // @[4_Mem.scala 70:27]
  reg [31:0] stageReg_csrAddr; // @[4_Mem.scala 70:27]
  reg [3:0] stageReg_excType; // @[4_Mem.scala 70:27]
  reg  stageReg_instState_commit; // @[4_Mem.scala 70:27]
  reg [31:0] stageReg_instState_pc; // @[4_Mem.scala 70:27]
  reg [31:0] stageReg_instState_inst; // @[4_Mem.scala 70:27]
  wire  _illgSret_T = stageReg_excType == 4'h3; // @[4_Mem.scala 82:38]
  wire  _illgSret_T_1 = io_csrMode == 2'h0; // @[4_Mem.scala 82:65]
  wire  illgSret = stageReg_excType == 4'h3 & io_csrMode == 2'h0; // @[4_Mem.scala 82:51]
  wire  _illgMret_T = stageReg_excType == 4'h4; // @[4_Mem.scala 83:38]
  wire  illgMret = stageReg_excType == 4'h4 & io_csrMode != 2'h3; // @[4_Mem.scala 83:51]
  wire  illgSpriv = stageReg_excType == 4'ha & _illgSret_T_1; // @[4_Mem.scala 84:52]
  wire  _instIllg_T_1 = stageReg_excType == 4'h5 | illgSret; // @[4_Mem.scala 87:52]
  wire  instIllg = _instIllg_T_1 | illgMret | illgSpriv; // @[4_Mem.scala 88:42]
  wire  _excOther_T_1 = stageReg_excType == 4'h2; // @[4_Mem.scala 90:38]
  wire  _excOther_T_2 = stageReg_excType == 4'h1 | _excOther_T_1; // @[4_Mem.scala 89:52]
  wire  _excOther_T_4 = _excOther_T_2 | _illgSret_T; // @[4_Mem.scala 90:51]
  wire  excOther = _excOther_T_4 | _illgMret_T; // @[4_Mem.scala 91:51]
  wire  hasTrap = (instIllg | excOther) & stageReg_instState_inst != 32'h0; // @[4_Mem.scala 93:44]
  wire [30:0] _cause_T_2 = io_csrMode == 2'h1 ? 31'h9 : 31'hb; // @[4_Mem.scala 98:32]
  wire [30:0] _cause_T_3 = _illgSret_T_1 ? 31'h8 : _cause_T_2; // @[4_Mem.scala 96:28]
  wire [30:0] _cause_T_5 = 4'h1 == stageReg_excType ? _cause_T_3 : 31'h0; // @[Mux.scala 81:58]
  wire [30:0] cause = 4'h2 == stageReg_excType ? 31'h3 : _cause_T_5; // @[Mux.scala 81:58]
  wire  _lsuSend_T = lsu_io_req_ready & lsu_io_req_valid; // @[Decoupled.scala 51:35]
  reg  lsuSend; // @[Reg.scala 35:20]
  wire  _GEN_48 = _lsuSend_T | lsuSend; // @[Reg.scala 36:18 35:20 36:22]
  LSU_1 lsu ( // @[4_Mem.scala 146:21]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_req_ready(lsu_io_req_ready),
    .io_req_valid(lsu_io_req_valid),
    .io_req_bits_addr(lsu_io_req_bits_addr),
    .io_req_bits_wdata(lsu_io_req_bits_wdata),
    .io_req_bits_lsuOp(lsu_io_req_bits_lsuOp),
    .io_resp_valid(lsu_io_resp_valid),
    .io_resp_bits_rdata(lsu_io_resp_bits_rdata),
    .io_cache_read_req_ready(lsu_io_cache_read_req_ready),
    .io_cache_read_req_valid(lsu_io_cache_read_req_valid),
    .io_cache_read_req_bits_addr(lsu_io_cache_read_req_bits_addr),
    .io_cache_read_resp_ready(lsu_io_cache_read_resp_ready),
    .io_cache_read_resp_valid(lsu_io_cache_read_resp_valid),
    .io_cache_read_resp_bits_data(lsu_io_cache_read_resp_bits_data),
    .io_cache_write_req_ready(lsu_io_cache_write_req_ready),
    .io_cache_write_req_valid(lsu_io_cache_write_req_valid),
    .io_cache_write_req_bits_addr(lsu_io_cache_write_req_bits_addr),
    .io_cache_write_req_bits_data(lsu_io_cache_write_req_bits_data),
    .io_cache_write_req_bits_mask(lsu_io_cache_write_req_bits_mask),
    .io_cache_write_resp_ready(lsu_io_cache_write_resp_ready),
    .io_cache_write_resp_valid(lsu_io_cache_write_resp_valid)
  );
  DCache dcache ( // @[4_Mem.scala 165:24]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_read_req_ready(dcache_io_read_req_ready),
    .io_read_req_valid(dcache_io_read_req_valid),
    .io_read_req_bits_addr(dcache_io_read_req_bits_addr),
    .io_read_resp_valid(dcache_io_read_resp_valid),
    .io_read_resp_bits_data(dcache_io_read_resp_bits_data),
    .io_write_req_ready(dcache_io_write_req_ready),
    .io_write_req_valid(dcache_io_write_req_valid),
    .io_write_req_bits_addr(dcache_io_write_req_bits_addr),
    .io_write_req_bits_data(dcache_io_write_req_bits_data),
    .io_write_req_bits_mask(dcache_io_write_req_bits_mask),
    .io_write_resp_valid(dcache_io_write_resp_valid),
    .io_tlbus_req_ready(dcache_io_tlbus_req_ready),
    .io_tlbus_req_valid(dcache_io_tlbus_req_valid),
    .io_tlbus_req_bits_opcode(dcache_io_tlbus_req_bits_opcode),
    .io_tlbus_req_bits_address(dcache_io_tlbus_req_bits_address),
    .io_tlbus_req_bits_data(dcache_io_tlbus_req_bits_data),
    .io_tlbus_resp_ready(dcache_io_tlbus_resp_ready),
    .io_tlbus_resp_valid(dcache_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(dcache_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(dcache_io_tlbus_resp_bits_data)
  );
  assign io_in_ready = ~stall & _io_in_ready_T_2; // @[4_Mem.scala 68:42]
  assign io_out_valid = ~stall; // @[4_Mem.scala 185:32]
  assign io_out_bits_resultSrc = stageReg_resultSrc; // @[4_Mem.scala 172:29]
  assign io_out_bits_regWrEn = stageReg_regWrEn; // @[4_Mem.scala 173:29]
  assign io_out_bits_aluOut = stageReg_aluOut; // @[4_Mem.scala 174:29]
  assign io_out_bits_pcNext4 = stageReg_pcNext4; // @[4_Mem.scala 175:29]
  assign io_out_bits_csrOp = stageReg_csrOp; // @[4_Mem.scala 115:29]
  assign io_out_bits_csrWrEn = stageReg_csrWrEn; // @[4_Mem.scala 116:29]
  assign io_out_bits_csrRdData = stageReg_csrRdData; // @[4_Mem.scala 117:29]
  assign io_out_bits_csrWrData = stageReg_csrWrData; // @[4_Mem.scala 118:29]
  assign io_out_bits_csrAddr = stageReg_csrAddr[11:0]; // @[4_Mem.scala 119:29]
  assign io_out_bits_instState_commit = stageReg_instState_commit; // @[4_Mem.scala 176:29]
  assign io_out_bits_instState_pc = stageReg_instState_pc; // @[4_Mem.scala 176:29]
  assign io_out_bits_instState_inst = stageReg_instState_inst; // @[4_Mem.scala 176:29]
  assign io_lsuData = lsu_io_resp_bits_rdata; // @[4_Mem.scala 163:29]
  assign io_lsuOK = lsu_io_resp_valid; // @[4_Mem.scala 162:29]
  assign io_tlbus_req_valid = dcache_io_tlbus_req_valid; // @[4_Mem.scala 168:21]
  assign io_tlbus_req_bits_opcode = dcache_io_tlbus_req_bits_opcode; // @[4_Mem.scala 168:21]
  assign io_tlbus_req_bits_address = dcache_io_tlbus_req_bits_address; // @[4_Mem.scala 168:21]
  assign io_tlbus_req_bits_data = dcache_io_tlbus_req_bits_data; // @[4_Mem.scala 168:21]
  assign io_hazard_rd = stageReg_instState_inst[11:7]; // @[util.scala 71:31]
  assign io_hazard_rdVal = stageReg_aluOut; // @[4_Mem.scala 183:29]
  assign io_hazard_regWrEn = stageReg_regWrEn; // @[4_Mem.scala 182:29]
  assign io_excp_valid = ~io_csrBusy & hasTrap & _io_in_ready_T; // @[4_Mem.scala 109:55]
  assign io_excp_bits_isMret = stageReg_excType == 4'h4; // @[4_Mem.scala 112:49]
  assign io_excp_bits_isSret = stageReg_excType == 4'h3; // @[4_Mem.scala 113:49]
  assign io_excp_bits_excCause = stageReg_csrWrEn & ~stageReg_csrValid ? 31'h2 : cause; // @[4_Mem.scala 105:35]
  assign io_excp_bits_excPc = stageReg_instState_pc; // @[4_Mem.scala 110:29]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_req_valid = stageReg_instState_commit & validLsuOp & ~lsuSend; // @[4_Mem.scala 157:72]
  assign lsu_io_req_bits_addr = stageReg_aluOut; // @[4_Mem.scala 158:29]
  assign lsu_io_req_bits_wdata = stageReg_data2; // @[4_Mem.scala 159:29]
  assign lsu_io_req_bits_lsuOp = stageReg_lsuOp; // @[4_Mem.scala 161:29]
  assign lsu_io_cache_read_req_ready = dcache_io_read_req_ready; // @[4_Mem.scala 166:23]
  assign lsu_io_cache_read_resp_valid = dcache_io_read_resp_valid; // @[4_Mem.scala 166:23]
  assign lsu_io_cache_read_resp_bits_data = dcache_io_read_resp_bits_data; // @[4_Mem.scala 166:23]
  assign lsu_io_cache_write_req_ready = dcache_io_write_req_ready; // @[4_Mem.scala 167:24]
  assign lsu_io_cache_write_resp_valid = dcache_io_write_resp_valid; // @[4_Mem.scala 167:24]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_read_req_valid = lsu_io_cache_read_req_valid; // @[4_Mem.scala 166:23]
  assign dcache_io_read_req_bits_addr = lsu_io_cache_read_req_bits_addr; // @[4_Mem.scala 166:23]
  assign dcache_io_write_req_valid = lsu_io_cache_write_req_valid; // @[4_Mem.scala 167:24]
  assign dcache_io_write_req_bits_addr = lsu_io_cache_write_req_bits_addr; // @[4_Mem.scala 167:24]
  assign dcache_io_write_req_bits_data = lsu_io_cache_write_req_bits_data; // @[4_Mem.scala 167:24]
  assign dcache_io_write_req_bits_mask = lsu_io_cache_write_req_bits_mask; // @[4_Mem.scala 167:24]
  assign dcache_io_tlbus_req_ready = io_tlbus_req_ready; // @[4_Mem.scala 168:21]
  assign dcache_io_tlbus_resp_valid = io_tlbus_resp_valid; // @[4_Mem.scala 168:21]
  assign dcache_io_tlbus_resp_bits_opcode = io_tlbus_resp_bits_opcode; // @[4_Mem.scala 168:21]
  assign dcache_io_tlbus_resp_bits_data = io_tlbus_resp_bits_data; // @[4_Mem.scala 168:21]
  always @(posedge clock) begin
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_lsuOp <= 5'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_lsuOp <= 5'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_lsuOp <= io_in_bits_lsuOp;
      end else begin
        stageReg_lsuOp <= 5'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_lsuOp <= 5'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_resultSrc <= 2'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_resultSrc <= 2'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_resultSrc <= io_in_bits_resultSrc;
      end else begin
        stageReg_resultSrc <= 2'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_resultSrc <= 2'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_regWrEn <= 1'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_regWrEn <= 1'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      stageReg_regWrEn <= io_in_bits_instState_commit & io_in_bits_regWrEn; // @[4_Mem.scala 72:18]
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_regWrEn <= 1'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_aluOut <= 32'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_aluOut <= 32'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_aluOut <= io_in_bits_aluOut;
      end else begin
        stageReg_aluOut <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_aluOut <= 32'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_data2 <= 32'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_data2 <= 32'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_data2 <= io_in_bits_data2;
      end else begin
        stageReg_data2 <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_data2 <= 32'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_pcNext4 <= 32'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_pcNext4 <= 32'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_pcNext4 <= io_in_bits_pcNext4;
      end else begin
        stageReg_pcNext4 <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_pcNext4 <= 32'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_csrOp <= 3'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_csrOp <= 3'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_csrOp <= io_in_bits_csrOp;
      end else begin
        stageReg_csrOp <= 3'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_csrOp <= 3'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_csrWrEn <= 1'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_csrWrEn <= 1'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      stageReg_csrWrEn <= io_in_bits_instState_commit & io_in_bits_csrWrEn; // @[4_Mem.scala 72:18]
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_csrWrEn <= 1'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_csrValid <= 1'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_csrValid <= 1'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      stageReg_csrValid <= io_in_bits_instState_commit & io_in_bits_csrValid; // @[4_Mem.scala 72:18]
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_csrValid <= 1'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_csrRdData <= 32'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_csrRdData <= 32'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_csrRdData <= io_in_bits_csrRdData;
      end else begin
        stageReg_csrRdData <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_csrRdData <= 32'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_csrWrData <= 32'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_csrWrData <= 32'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_csrWrData <= io_in_bits_csrWrData;
      end else begin
        stageReg_csrWrData <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_csrWrData <= 32'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_csrAddr <= 32'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_csrAddr <= 32'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_csrAddr <= io_in_bits_csrAddr;
      end else begin
        stageReg_csrAddr <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_csrAddr <= 32'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_excType <= 4'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_excType <= 4'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_excType <= io_in_bits_excType;
      end else begin
        stageReg_excType <= 4'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_excType <= 4'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_instState_commit <= 1'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_instState_commit <= 1'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      stageReg_instState_commit <= io_in_bits_instState_commit; // @[4_Mem.scala 72:18]
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_instState_commit <= 1'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_instState_pc <= 32'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_instState_pc <= 32'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_instState_pc <= io_in_bits_instState_pc;
      end else begin
        stageReg_instState_pc <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_instState_pc <= 32'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[4_Mem.scala 70:27]
      stageReg_instState_inst <= 32'h0; // @[4_Mem.scala 70:27]
    end else if (io_ctrl_flush & _io_in_ready_T) begin // @[4_Mem.scala 77:27]
      stageReg_instState_inst <= 32'h0; // @[4_Mem.scala 77:38]
    end else if (io_in_ready) begin // @[4_Mem.scala 71:23]
      if (io_in_bits_instState_commit) begin // @[4_Mem.scala 72:24]
        stageReg_instState_inst <= io_in_bits_instState_inst;
      end else begin
        stageReg_instState_inst <= 32'h0;
      end
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 73:28]
      stageReg_instState_inst <= 32'h0; // @[4_Mem.scala 74:18]
    end
    if (reset) begin // @[Reg.scala 35:20]
      lsuSend <= 1'h0; // @[Reg.scala 35:20]
    end else if (_io_in_ready_T_2) begin // @[4_Mem.scala 156:23]
      lsuSend <= 1'h0; // @[4_Mem.scala 156:33]
    end else begin
      lsuSend <= _GEN_48;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stageReg_lsuOp = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  stageReg_resultSrc = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  stageReg_regWrEn = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  stageReg_aluOut = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  stageReg_data2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  stageReg_pcNext4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  stageReg_csrOp = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  stageReg_csrWrEn = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  stageReg_csrValid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  stageReg_csrRdData = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  stageReg_csrWrData = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  stageReg_csrAddr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  stageReg_excType = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  stageReg_instState_commit = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  stageReg_instState_pc = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  stageReg_instState_inst = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  lsuSend = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteBack(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [1:0]  io_in_bits_resultSrc,
  input         io_in_bits_regWrEn,
  input  [31:0] io_in_bits_aluOut,
  input  [31:0] io_in_bits_pcNext4,
  input  [2:0]  io_in_bits_csrOp,
  input         io_in_bits_csrWrEn,
  input  [31:0] io_in_bits_csrRdData,
  input  [31:0] io_in_bits_csrWrData,
  input  [11:0] io_in_bits_csrAddr,
  input         io_in_bits_instState_commit,
  input  [31:0] io_in_bits_instState_pc,
  input  [31:0] io_in_bits_instState_inst,
  output        io_instState_commit,
  output [31:0] io_instState_pc,
  output [31:0] io_instState_inst,
  output [4:0]  io_hazard_rd,
  output [31:0] io_hazard_rdVal,
  output        io_hazard_regWrEn,
  output [4:0]  io_regfile_rd,
  output        io_regfile_regWrEn,
  output [31:0] io_regfile_regWrData,
  output [2:0]  io_csrWrite_op,
  output [11:0] io_csrWrite_addr,
  output [31:0] io_csrWrite_data,
  output        io_csrWrite_retired,
  input  [31:0] io_lsuData
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  writebackLatch = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  reg [1:0] stageReg_resultSrc; // @[5_WriteBack.scala 44:27]
  reg  stageReg_regWrEn; // @[5_WriteBack.scala 44:27]
  reg [31:0] stageReg_aluOut; // @[5_WriteBack.scala 44:27]
  reg [31:0] stageReg_pcNext4; // @[5_WriteBack.scala 44:27]
  reg [2:0] stageReg_csrOp; // @[5_WriteBack.scala 44:27]
  reg  stageReg_csrWrEn; // @[5_WriteBack.scala 44:27]
  reg [31:0] stageReg_csrRdData; // @[5_WriteBack.scala 44:27]
  reg [31:0] stageReg_csrWrData; // @[5_WriteBack.scala 44:27]
  reg [11:0] stageReg_csrAddr; // @[5_WriteBack.scala 44:27]
  reg  stageReg_instState_commit; // @[5_WriteBack.scala 44:27]
  reg [31:0] stageReg_instState_pc; // @[5_WriteBack.scala 44:27]
  reg [31:0] stageReg_instState_inst; // @[5_WriteBack.scala 44:27]
  wire  _GEN_13 = writebackLatch & (io_in_bits_instState_commit & io_in_bits_regWrEn); // @[5_WriteBack.scala 45:26 46:18]
  wire  _GEN_17 = writebackLatch & (io_in_bits_instState_commit & io_in_bits_csrWrEn); // @[5_WriteBack.scala 45:26 46:18]
  wire  _GEN_21 = writebackLatch & io_in_bits_instState_commit; // @[5_WriteBack.scala 45:26 46:18]
  wire [31:0] _rdVal_T_1 = 2'h1 == stageReg_resultSrc ? io_lsuData : stageReg_aluOut; // @[Mux.scala 81:58]
  wire [31:0] _rdVal_T_3 = 2'h2 == stageReg_resultSrc ? stageReg_pcNext4 : _rdVal_T_1; // @[Mux.scala 81:58]
  assign io_in_ready = io_in_valid; // @[5_WriteBack.scala 42:27]
  assign io_instState_commit = stageReg_instState_commit; // @[5_WriteBack.scala 73:55]
  assign io_instState_pc = stageReg_instState_pc; // @[5_WriteBack.scala 72:26]
  assign io_instState_inst = stageReg_instState_inst; // @[5_WriteBack.scala 72:26]
  assign io_hazard_rd = stageReg_instState_inst[11:7]; // @[util.scala 71:31]
  assign io_hazard_rdVal = 2'h3 == stageReg_resultSrc ? stageReg_csrRdData : _rdVal_T_3; // @[Mux.scala 81:58]
  assign io_hazard_regWrEn = stageReg_regWrEn; // @[5_WriteBack.scala 78:26]
  assign io_regfile_rd = stageReg_instState_inst[11:7]; // @[util.scala 71:31]
  assign io_regfile_regWrEn = stageReg_regWrEn & stageReg_instState_commit; // @[5_WriteBack.scala 64:46]
  assign io_regfile_regWrData = 2'h3 == stageReg_resultSrc ? stageReg_csrRdData : _rdVal_T_3; // @[Mux.scala 81:58]
  assign io_csrWrite_op = stageReg_csrWrEn ? stageReg_csrOp : 3'h1; // @[5_WriteBack.scala 69:32]
  assign io_csrWrite_addr = stageReg_csrAddr; // @[5_WriteBack.scala 67:26]
  assign io_csrWrite_data = stageReg_csrWrData; // @[5_WriteBack.scala 68:26]
  assign io_csrWrite_retired = stageReg_instState_commit; // @[5_WriteBack.scala 70:55]
  always @(posedge clock) begin
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_resultSrc <= 2'h0; // @[5_WriteBack.scala 44:27]
    end else if (writebackLatch) begin // @[5_WriteBack.scala 45:26]
      if (io_in_bits_instState_commit) begin // @[5_WriteBack.scala 46:24]
        stageReg_resultSrc <= io_in_bits_resultSrc;
      end else begin
        stageReg_resultSrc <= 2'h0;
      end
    end else begin
      stageReg_resultSrc <= 2'h0;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_regWrEn <= 1'h0; // @[5_WriteBack.scala 44:27]
    end else begin
      stageReg_regWrEn <= _GEN_13;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_aluOut <= 32'h0; // @[5_WriteBack.scala 44:27]
    end else if (writebackLatch) begin // @[5_WriteBack.scala 45:26]
      if (io_in_bits_instState_commit) begin // @[5_WriteBack.scala 46:24]
        stageReg_aluOut <= io_in_bits_aluOut;
      end else begin
        stageReg_aluOut <= 32'h0;
      end
    end else begin
      stageReg_aluOut <= 32'h0;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_pcNext4 <= 32'h0; // @[5_WriteBack.scala 44:27]
    end else if (writebackLatch) begin // @[5_WriteBack.scala 45:26]
      if (io_in_bits_instState_commit) begin // @[5_WriteBack.scala 46:24]
        stageReg_pcNext4 <= io_in_bits_pcNext4;
      end else begin
        stageReg_pcNext4 <= 32'h0;
      end
    end else begin
      stageReg_pcNext4 <= 32'h0;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_csrOp <= 3'h0; // @[5_WriteBack.scala 44:27]
    end else if (writebackLatch) begin // @[5_WriteBack.scala 45:26]
      if (io_in_bits_instState_commit) begin // @[5_WriteBack.scala 46:24]
        stageReg_csrOp <= io_in_bits_csrOp;
      end else begin
        stageReg_csrOp <= 3'h0;
      end
    end else begin
      stageReg_csrOp <= 3'h0;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_csrWrEn <= 1'h0; // @[5_WriteBack.scala 44:27]
    end else begin
      stageReg_csrWrEn <= _GEN_17;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_csrRdData <= 32'h0; // @[5_WriteBack.scala 44:27]
    end else if (writebackLatch) begin // @[5_WriteBack.scala 45:26]
      if (io_in_bits_instState_commit) begin // @[5_WriteBack.scala 46:24]
        stageReg_csrRdData <= io_in_bits_csrRdData;
      end else begin
        stageReg_csrRdData <= 32'h0;
      end
    end else begin
      stageReg_csrRdData <= 32'h0;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_csrWrData <= 32'h0; // @[5_WriteBack.scala 44:27]
    end else if (writebackLatch) begin // @[5_WriteBack.scala 45:26]
      if (io_in_bits_instState_commit) begin // @[5_WriteBack.scala 46:24]
        stageReg_csrWrData <= io_in_bits_csrWrData;
      end else begin
        stageReg_csrWrData <= 32'h0;
      end
    end else begin
      stageReg_csrWrData <= 32'h0;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_csrAddr <= 12'h0; // @[5_WriteBack.scala 44:27]
    end else if (writebackLatch) begin // @[5_WriteBack.scala 45:26]
      if (io_in_bits_instState_commit) begin // @[5_WriteBack.scala 46:24]
        stageReg_csrAddr <= io_in_bits_csrAddr;
      end else begin
        stageReg_csrAddr <= 12'h0;
      end
    end else begin
      stageReg_csrAddr <= 12'h0;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_instState_commit <= 1'h0; // @[5_WriteBack.scala 44:27]
    end else begin
      stageReg_instState_commit <= _GEN_21;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_instState_pc <= 32'h0; // @[5_WriteBack.scala 44:27]
    end else if (writebackLatch) begin // @[5_WriteBack.scala 45:26]
      if (io_in_bits_instState_commit) begin // @[5_WriteBack.scala 46:24]
        stageReg_instState_pc <= io_in_bits_instState_pc;
      end else begin
        stageReg_instState_pc <= 32'h0;
      end
    end else begin
      stageReg_instState_pc <= 32'h0;
    end
    if (reset) begin // @[5_WriteBack.scala 44:27]
      stageReg_instState_inst <= 32'h0; // @[5_WriteBack.scala 44:27]
    end else if (writebackLatch) begin // @[5_WriteBack.scala 45:26]
      if (io_in_bits_instState_commit) begin // @[5_WriteBack.scala 46:24]
        stageReg_instState_inst <= io_in_bits_instState_inst;
      end else begin
        stageReg_instState_inst <= 32'h0;
      end
    end else begin
      stageReg_instState_inst <= 32'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stageReg_resultSrc = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  stageReg_regWrEn = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  stageReg_aluOut = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  stageReg_pcNext4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  stageReg_csrOp = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  stageReg_csrWrEn = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  stageReg_csrRdData = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  stageReg_csrWrData = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  stageReg_csrAddr = _RAND_8[11:0];
  _RAND_9 = {1{`RANDOM}};
  stageReg_instState_commit = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  stageReg_instState_pc = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  stageReg_instState_inst = _RAND_11[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineCtrl(
  input   io_in_brTaken,
  input   io_in_excpValid,
  output  io_out_decode_flush,
  output  io_out_execute_flush,
  output  io_out_memory_flush
);
  assign io_out_decode_flush = io_in_brTaken | io_in_excpValid; // @[PipelineCtrl.scala 35:38]
  assign io_out_execute_flush = io_in_excpValid; // @[PipelineCtrl.scala 36:26]
  assign io_out_memory_flush = io_in_excpValid; // @[PipelineCtrl.scala 37:25]
endmodule
module HazardUnit(
  input  [4:0]  io_in_decode_rs1,
  input  [4:0]  io_in_decode_rs2,
  input  [4:0]  io_in_execute_rs1,
  input  [4:0]  io_in_execute_rs2,
  input  [1:0]  io_in_execute_resultSrc,
  input  [4:0]  io_in_execute_rd,
  input  [4:0]  io_in_memory_rd,
  input  [31:0] io_in_memory_rdVal,
  input         io_in_memory_regWrEn,
  input  [4:0]  io_in_writeback_rd,
  input  [31:0] io_in_writeback_rdVal,
  input         io_in_writeback_regWrEn,
  output [1:0]  io_out_execute_aluSrc1,
  output [1:0]  io_out_execute_aluSrc2,
  output [31:0] io_out_execute_rdValM,
  output [31:0] io_out_execute_rdValW,
  output        io_out_decode_stall
);
  wire  _fwMem2ExeRs1_T_2 = io_in_memory_rd != 5'h0; // @[HazardUnit.scala 41:58]
  wire  fwMem2ExeRs1 = io_in_execute_rs1 == io_in_memory_rd & io_in_memory_regWrEn & io_in_memory_rd != 5'h0; // @[HazardUnit.scala 41:51]
  wire  fwMem2ExeRs2 = io_in_execute_rs2 == io_in_memory_rd & io_in_memory_regWrEn & _fwMem2ExeRs1_T_2; // @[HazardUnit.scala 43:51]
  wire  _fwWb2ExeRs1_T_2 = io_in_writeback_rd != 5'h0; // @[HazardUnit.scala 46:57]
  wire  fwWb2ExeRs1 = io_in_execute_rs1 == io_in_writeback_rd & io_in_writeback_regWrEn & io_in_writeback_rd != 5'h0; // @[HazardUnit.scala 46:50]
  wire  fwWb2ExeRs2 = io_in_execute_rs2 == io_in_writeback_rd & io_in_writeback_regWrEn & _fwWb2ExeRs1_T_2; // @[HazardUnit.scala 48:50]
  wire [1:0] _GEN_0 = fwWb2ExeRs1 ? 2'h2 : 2'h0; // @[HazardUnit.scala 54:25 51:28 55:32]
  wire [1:0] _GEN_1 = fwWb2ExeRs2 ? 2'h2 : 2'h0; // @[HazardUnit.scala 57:25 52:28 58:32]
  wire  _T_5 = io_in_execute_rd == io_in_decode_rs1 | io_in_execute_rd == io_in_decode_rs2; // @[HazardUnit.scala 79:27]
  assign io_out_execute_aluSrc1 = fwMem2ExeRs1 ? 2'h1 : _GEN_0; // @[HazardUnit.scala 62:26 63:32]
  assign io_out_execute_aluSrc2 = fwMem2ExeRs2 ? 2'h1 : _GEN_1; // @[HazardUnit.scala 65:26 66:32]
  assign io_out_execute_rdValM = io_in_memory_rdVal; // @[HazardUnit.scala 69:27]
  assign io_out_execute_rdValW = io_in_writeback_rdVal; // @[HazardUnit.scala 70:27]
  assign io_out_decode_stall = io_in_execute_resultSrc == 2'h1 & io_in_execute_rd != 5'h0 & _T_5; // @[HazardUnit.scala 77:25 78:51]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_r_0_addr,
  output [31:0] io_r_0_data,
  input  [4:0]  io_r_1_addr,
  output [31:0] io_r_1_data,
  input  [4:0]  io_w_0_addr,
  input         io_w_0_en,
  input  [31:0] io_w_0_data,
  output [31:0] regState_0_regState_0,
  output [31:0] regState_0_regState_1,
  output [31:0] regState_0_regState_2,
  output [31:0] regState_0_regState_3,
  output [31:0] regState_0_regState_4,
  output [31:0] regState_0_regState_5,
  output [31:0] regState_0_regState_6,
  output [31:0] regState_0_regState_7,
  output [31:0] regState_0_regState_8,
  output [31:0] regState_0_regState_9,
  output [31:0] regState_0_regState_10,
  output [31:0] regState_0_regState_11,
  output [31:0] regState_0_regState_12,
  output [31:0] regState_0_regState_13,
  output [31:0] regState_0_regState_14,
  output [31:0] regState_0_regState_15,
  output [31:0] regState_0_regState_16,
  output [31:0] regState_0_regState_17,
  output [31:0] regState_0_regState_18,
  output [31:0] regState_0_regState_19,
  output [31:0] regState_0_regState_20,
  output [31:0] regState_0_regState_21,
  output [31:0] regState_0_regState_22,
  output [31:0] regState_0_regState_23,
  output [31:0] regState_0_regState_24,
  output [31:0] regState_0_regState_25,
  output [31:0] regState_0_regState_26,
  output [31:0] regState_0_regState_27,
  output [31:0] regState_0_regState_28,
  output [31:0] regState_0_regState_29,
  output [31:0] regState_0_regState_30,
  output [31:0] regState_0_regState_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[RegFile.scala 31:17]
  reg [31:0] regs_1; // @[RegFile.scala 31:17]
  reg [31:0] regs_2; // @[RegFile.scala 31:17]
  reg [31:0] regs_3; // @[RegFile.scala 31:17]
  reg [31:0] regs_4; // @[RegFile.scala 31:17]
  reg [31:0] regs_5; // @[RegFile.scala 31:17]
  reg [31:0] regs_6; // @[RegFile.scala 31:17]
  reg [31:0] regs_7; // @[RegFile.scala 31:17]
  reg [31:0] regs_8; // @[RegFile.scala 31:17]
  reg [31:0] regs_9; // @[RegFile.scala 31:17]
  reg [31:0] regs_10; // @[RegFile.scala 31:17]
  reg [31:0] regs_11; // @[RegFile.scala 31:17]
  reg [31:0] regs_12; // @[RegFile.scala 31:17]
  reg [31:0] regs_13; // @[RegFile.scala 31:17]
  reg [31:0] regs_14; // @[RegFile.scala 31:17]
  reg [31:0] regs_15; // @[RegFile.scala 31:17]
  reg [31:0] regs_16; // @[RegFile.scala 31:17]
  reg [31:0] regs_17; // @[RegFile.scala 31:17]
  reg [31:0] regs_18; // @[RegFile.scala 31:17]
  reg [31:0] regs_19; // @[RegFile.scala 31:17]
  reg [31:0] regs_20; // @[RegFile.scala 31:17]
  reg [31:0] regs_21; // @[RegFile.scala 31:17]
  reg [31:0] regs_22; // @[RegFile.scala 31:17]
  reg [31:0] regs_23; // @[RegFile.scala 31:17]
  reg [31:0] regs_24; // @[RegFile.scala 31:17]
  reg [31:0] regs_25; // @[RegFile.scala 31:17]
  reg [31:0] regs_26; // @[RegFile.scala 31:17]
  reg [31:0] regs_27; // @[RegFile.scala 31:17]
  reg [31:0] regs_28; // @[RegFile.scala 31:17]
  reg [31:0] regs_29; // @[RegFile.scala 31:17]
  reg [31:0] regs_30; // @[RegFile.scala 31:17]
  reg [31:0] regs_31; // @[RegFile.scala 31:17]
  wire [31:0] _GEN_1 = reset ? 32'h0 : regs_1; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_2 = reset ? 32'h0 : regs_2; // @[RegFile.scala 32:22 37:11 31:17]
  wire [31:0] _GEN_3 = reset ? 32'h0 : regs_3; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_4 = reset ? 32'h0 : regs_4; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_5 = reset ? 32'h0 : regs_5; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_6 = reset ? 32'h0 : regs_6; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_7 = reset ? 32'h0 : regs_7; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_8 = reset ? 32'h0 : regs_8; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_9 = reset ? 32'h0 : regs_9; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_10 = reset ? 32'h0 : regs_10; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_11 = reset ? 32'h0 : regs_11; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_12 = reset ? 32'h0 : regs_12; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_13 = reset ? 32'h0 : regs_13; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_14 = reset ? 32'h0 : regs_14; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_15 = reset ? 32'h0 : regs_15; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_16 = reset ? 32'h0 : regs_16; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_17 = reset ? 32'h0 : regs_17; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_18 = reset ? 32'h0 : regs_18; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_19 = reset ? 32'h0 : regs_19; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_20 = reset ? 32'h0 : regs_20; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_21 = reset ? 32'h0 : regs_21; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_22 = reset ? 32'h0 : regs_22; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_23 = reset ? 32'h0 : regs_23; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_24 = reset ? 32'h0 : regs_24; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_25 = reset ? 32'h0 : regs_25; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_26 = reset ? 32'h0 : regs_26; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_27 = reset ? 32'h0 : regs_27; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_28 = reset ? 32'h0 : regs_28; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_29 = reset ? 32'h0 : regs_29; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_30 = reset ? 32'h0 : regs_30; // @[RegFile.scala 31:17 32:22 34:9]
  wire [31:0] _GEN_31 = reset ? 32'h0 : regs_31; // @[RegFile.scala 31:17 32:22 34:9]
  wire  _writeBypassVec_T_2 = io_w_0_addr != 5'h0; // @[RegFile.scala 45:67]
  wire  writeBypassVec_0 = io_w_0_en & io_r_0_addr == io_w_0_addr & io_w_0_addr != 5'h0; // @[RegFile.scala 45:51]
  wire  writeBypassVec_1 = io_w_0_en & io_r_1_addr == io_w_0_addr & io_w_0_addr != 5'h0; // @[RegFile.scala 45:51]
  wire [31:0] _GEN_32 = regs_0; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_33 = 5'h1 == io_r_0_addr ? regs_1 : regs_0; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_34 = 5'h2 == io_r_0_addr ? regs_2 : _GEN_33; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_35 = 5'h3 == io_r_0_addr ? regs_3 : _GEN_34; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_36 = 5'h4 == io_r_0_addr ? regs_4 : _GEN_35; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_37 = 5'h5 == io_r_0_addr ? regs_5 : _GEN_36; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_38 = 5'h6 == io_r_0_addr ? regs_6 : _GEN_37; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_39 = 5'h7 == io_r_0_addr ? regs_7 : _GEN_38; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_40 = 5'h8 == io_r_0_addr ? regs_8 : _GEN_39; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_41 = 5'h9 == io_r_0_addr ? regs_9 : _GEN_40; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_42 = 5'ha == io_r_0_addr ? regs_10 : _GEN_41; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_43 = 5'hb == io_r_0_addr ? regs_11 : _GEN_42; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_44 = 5'hc == io_r_0_addr ? regs_12 : _GEN_43; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_45 = 5'hd == io_r_0_addr ? regs_13 : _GEN_44; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_46 = 5'he == io_r_0_addr ? regs_14 : _GEN_45; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_47 = 5'hf == io_r_0_addr ? regs_15 : _GEN_46; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_48 = 5'h10 == io_r_0_addr ? regs_16 : _GEN_47; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_49 = 5'h11 == io_r_0_addr ? regs_17 : _GEN_48; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_50 = 5'h12 == io_r_0_addr ? regs_18 : _GEN_49; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_51 = 5'h13 == io_r_0_addr ? regs_19 : _GEN_50; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_52 = 5'h14 == io_r_0_addr ? regs_20 : _GEN_51; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_53 = 5'h15 == io_r_0_addr ? regs_21 : _GEN_52; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_54 = 5'h16 == io_r_0_addr ? regs_22 : _GEN_53; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_55 = 5'h17 == io_r_0_addr ? regs_23 : _GEN_54; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_56 = 5'h18 == io_r_0_addr ? regs_24 : _GEN_55; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_57 = 5'h19 == io_r_0_addr ? regs_25 : _GEN_56; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_58 = 5'h1a == io_r_0_addr ? regs_26 : _GEN_57; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_59 = 5'h1b == io_r_0_addr ? regs_27 : _GEN_58; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_60 = 5'h1c == io_r_0_addr ? regs_28 : _GEN_59; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_61 = 5'h1d == io_r_0_addr ? regs_29 : _GEN_60; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_62 = 5'h1e == io_r_0_addr ? regs_30 : _GEN_61; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_63 = 5'h1f == io_r_0_addr ? regs_31 : _GEN_62; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_67 = 5'h1 == io_r_1_addr ? regs_1 : regs_0; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_68 = 5'h2 == io_r_1_addr ? regs_2 : _GEN_67; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_69 = 5'h3 == io_r_1_addr ? regs_3 : _GEN_68; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_70 = 5'h4 == io_r_1_addr ? regs_4 : _GEN_69; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_71 = 5'h5 == io_r_1_addr ? regs_5 : _GEN_70; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_72 = 5'h6 == io_r_1_addr ? regs_6 : _GEN_71; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_73 = 5'h7 == io_r_1_addr ? regs_7 : _GEN_72; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_74 = 5'h8 == io_r_1_addr ? regs_8 : _GEN_73; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_75 = 5'h9 == io_r_1_addr ? regs_9 : _GEN_74; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_76 = 5'ha == io_r_1_addr ? regs_10 : _GEN_75; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_77 = 5'hb == io_r_1_addr ? regs_11 : _GEN_76; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_78 = 5'hc == io_r_1_addr ? regs_12 : _GEN_77; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_79 = 5'hd == io_r_1_addr ? regs_13 : _GEN_78; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_80 = 5'he == io_r_1_addr ? regs_14 : _GEN_79; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_81 = 5'hf == io_r_1_addr ? regs_15 : _GEN_80; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_82 = 5'h10 == io_r_1_addr ? regs_16 : _GEN_81; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_83 = 5'h11 == io_r_1_addr ? regs_17 : _GEN_82; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_84 = 5'h12 == io_r_1_addr ? regs_18 : _GEN_83; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_85 = 5'h13 == io_r_1_addr ? regs_19 : _GEN_84; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_86 = 5'h14 == io_r_1_addr ? regs_20 : _GEN_85; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_87 = 5'h15 == io_r_1_addr ? regs_21 : _GEN_86; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_88 = 5'h16 == io_r_1_addr ? regs_22 : _GEN_87; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_89 = 5'h17 == io_r_1_addr ? regs_23 : _GEN_88; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_90 = 5'h18 == io_r_1_addr ? regs_24 : _GEN_89; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_91 = 5'h19 == io_r_1_addr ? regs_25 : _GEN_90; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_92 = 5'h1a == io_r_1_addr ? regs_26 : _GEN_91; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_93 = 5'h1b == io_r_1_addr ? regs_27 : _GEN_92; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_94 = 5'h1c == io_r_1_addr ? regs_28 : _GEN_93; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_95 = 5'h1d == io_r_1_addr ? regs_29 : _GEN_94; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_96 = 5'h1e == io_r_1_addr ? regs_30 : _GEN_95; // @[RegFile.scala 53:{22,22}]
  wire [31:0] _GEN_97 = 5'h1f == io_r_1_addr ? regs_31 : _GEN_96; // @[RegFile.scala 53:{22,22}]
  wire [31:0] regState_regState_0 = regs_0; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_1 = regs_1; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_2 = regs_2; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_3 = regs_3; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_4 = regs_4; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_5 = regs_5; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_6 = regs_6; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_7 = regs_7; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_8 = regs_8; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_9 = regs_9; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_10 = regs_10; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_11 = regs_11; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_12 = regs_12; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_13 = regs_13; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_14 = regs_14; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_15 = regs_15; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_16 = regs_16; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_17 = regs_17; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_18 = regs_18; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_19 = regs_19; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_20 = regs_20; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_21 = regs_21; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_22 = regs_22; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_23 = regs_23; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_24 = regs_24; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_25 = regs_25; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_26 = regs_26; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_27 = regs_27; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_28 = regs_28; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_29 = regs_29; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_30 = regs_30; // @[RegFile.scala 108:24 110:9]
  wire [31:0] regState_regState_31 = regs_31; // @[RegFile.scala 108:24 110:9]
  assign io_r_0_data = writeBypassVec_0 ? io_w_0_data : _GEN_63; // @[RegFile.scala 50:31 51:22 53:22]
  assign io_r_1_data = writeBypassVec_1 ? io_w_0_data : _GEN_97; // @[RegFile.scala 50:31 51:22 53:22]
  assign regState_0_regState_0 = _GEN_32;
  assign regState_0_regState_1 = regState_regState_1;
  assign regState_0_regState_2 = regState_regState_2;
  assign regState_0_regState_3 = regState_regState_3;
  assign regState_0_regState_4 = regState_regState_4;
  assign regState_0_regState_5 = regState_regState_5;
  assign regState_0_regState_6 = regState_regState_6;
  assign regState_0_regState_7 = regState_regState_7;
  assign regState_0_regState_8 = regState_regState_8;
  assign regState_0_regState_9 = regState_regState_9;
  assign regState_0_regState_10 = regState_regState_10;
  assign regState_0_regState_11 = regState_regState_11;
  assign regState_0_regState_12 = regState_regState_12;
  assign regState_0_regState_13 = regState_regState_13;
  assign regState_0_regState_14 = regState_regState_14;
  assign regState_0_regState_15 = regState_regState_15;
  assign regState_0_regState_16 = regState_regState_16;
  assign regState_0_regState_17 = regState_regState_17;
  assign regState_0_regState_18 = regState_regState_18;
  assign regState_0_regState_19 = regState_regState_19;
  assign regState_0_regState_20 = regState_regState_20;
  assign regState_0_regState_21 = regState_regState_21;
  assign regState_0_regState_22 = regState_regState_22;
  assign regState_0_regState_23 = regState_regState_23;
  assign regState_0_regState_24 = regState_regState_24;
  assign regState_0_regState_25 = regState_regState_25;
  assign regState_0_regState_26 = regState_regState_26;
  assign regState_0_regState_27 = regState_regState_27;
  assign regState_0_regState_28 = regState_regState_28;
  assign regState_0_regState_29 = regState_regState_29;
  assign regState_0_regState_30 = regState_regState_30;
  assign regState_0_regState_31 = regState_regState_31;
  always @(posedge clock) begin
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h0 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_0 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_0 <= 32'h0; // @[RegFile.scala 40:11]
      end
    end else begin
      regs_0 <= 32'h0; // @[RegFile.scala 40:11]
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h1 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_1 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_1 <= _GEN_1;
      end
    end else begin
      regs_1 <= _GEN_1;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h2 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_2 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_2 <= _GEN_2;
      end
    end else begin
      regs_2 <= _GEN_2;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h3 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_3 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_3 <= _GEN_3;
      end
    end else begin
      regs_3 <= _GEN_3;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h4 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_4 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_4 <= _GEN_4;
      end
    end else begin
      regs_4 <= _GEN_4;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h5 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_5 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_5 <= _GEN_5;
      end
    end else begin
      regs_5 <= _GEN_5;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h6 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_6 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_6 <= _GEN_6;
      end
    end else begin
      regs_6 <= _GEN_6;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h7 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_7 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_7 <= _GEN_7;
      end
    end else begin
      regs_7 <= _GEN_7;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h8 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_8 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_8 <= _GEN_8;
      end
    end else begin
      regs_8 <= _GEN_8;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h9 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_9 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_9 <= _GEN_9;
      end
    end else begin
      regs_9 <= _GEN_9;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'ha == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_10 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_10 <= _GEN_10;
      end
    end else begin
      regs_10 <= _GEN_10;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'hb == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_11 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_11 <= _GEN_11;
      end
    end else begin
      regs_11 <= _GEN_11;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'hc == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_12 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_12 <= _GEN_12;
      end
    end else begin
      regs_12 <= _GEN_12;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'hd == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_13 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_13 <= _GEN_13;
      end
    end else begin
      regs_13 <= _GEN_13;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'he == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_14 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_14 <= _GEN_14;
      end
    end else begin
      regs_14 <= _GEN_14;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'hf == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_15 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_15 <= _GEN_15;
      end
    end else begin
      regs_15 <= _GEN_15;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h10 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_16 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_16 <= _GEN_16;
      end
    end else begin
      regs_16 <= _GEN_16;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h11 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_17 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_17 <= _GEN_17;
      end
    end else begin
      regs_17 <= _GEN_17;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h12 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_18 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_18 <= _GEN_18;
      end
    end else begin
      regs_18 <= _GEN_18;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h13 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_19 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_19 <= _GEN_19;
      end
    end else begin
      regs_19 <= _GEN_19;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h14 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_20 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_20 <= _GEN_20;
      end
    end else begin
      regs_20 <= _GEN_20;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h15 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_21 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_21 <= _GEN_21;
      end
    end else begin
      regs_21 <= _GEN_21;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h16 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_22 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_22 <= _GEN_22;
      end
    end else begin
      regs_22 <= _GEN_22;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h17 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_23 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_23 <= _GEN_23;
      end
    end else begin
      regs_23 <= _GEN_23;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h18 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_24 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_24 <= _GEN_24;
      end
    end else begin
      regs_24 <= _GEN_24;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h19 == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_25 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_25 <= _GEN_25;
      end
    end else begin
      regs_25 <= _GEN_25;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h1a == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_26 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_26 <= _GEN_26;
      end
    end else begin
      regs_26 <= _GEN_26;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h1b == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_27 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_27 <= _GEN_27;
      end
    end else begin
      regs_27 <= _GEN_27;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h1c == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_28 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_28 <= _GEN_28;
      end
    end else begin
      regs_28 <= _GEN_28;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h1d == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_29 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_29 <= _GEN_29;
      end
    end else begin
      regs_29 <= _GEN_29;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h1e == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_30 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_30 <= _GEN_30;
      end
    end else begin
      regs_30 <= _GEN_30;
    end
    if (io_w_0_en & _writeBypassVec_T_2) begin // @[RegFile.scala 60:44]
      if (5'h1f == io_w_0_addr) begin // @[RegFile.scala 61:24]
        regs_31 <= io_w_0_data; // @[RegFile.scala 61:24]
      end else begin
        regs_31 <= _GEN_31;
      end
    end else begin
      regs_31 <= _GEN_31;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(regs_0 == 32'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed: zero reg must be 0 !\n    at RegFile.scala:41 assert(regs(0).asUInt === 0.U, \"zero reg must be 0 !\")\n"
            ); // @[RegFile.scala 41:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(regs_0 == 32'h0) & ~reset) begin
          $fatal; // @[RegFile.scala 41:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CsrFile(
  input         clock,
  input         reset,
  input  [2:0]  io_read_op,
  output        io_read_valid,
  input  [11:0] io_read_addr,
  output [31:0] io_read_data,
  input  [2:0]  io_write_op,
  input  [11:0] io_write_addr,
  input  [31:0] io_write_data,
  input         io_write_retired,
  input         io_except_valid,
  input         io_except_bits_isMret,
  input         io_except_bits_isSret,
  input  [30:0] io_except_bits_excCause,
  input  [31:0] io_except_bits_excPc,
  input  [31:0] io_except_bits_excValue,
  output [1:0]  io_mode,
  output        io_busy,
  output [31:0] io_mepc,
  output [31:0] io_trapVec,
  output [31:0] csrState_0_mcycle,
  output [31:0] csrState_0_mcycleh
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg  mcause_int; // @[CsrFile.scala 69:28]
  reg [30:0] mcause_code; // @[CsrFile.scala 69:28]
  reg  mstatus_sum; // @[CsrFile.scala 70:28]
  reg [1:0] mstatus_mpp; // @[CsrFile.scala 70:28]
  reg  mstatus_spp; // @[CsrFile.scala 70:28]
  reg  mstatus_mpie; // @[CsrFile.scala 70:28]
  reg  mstatus_spie; // @[CsrFile.scala 70:28]
  reg  mstatus_mie; // @[CsrFile.scala 70:28]
  reg  mstatus_sie; // @[CsrFile.scala 70:28]
  reg [29:0] mtvec_base; // @[CsrFile.scala 71:28]
  reg [1:0] mtvec_mode; // @[CsrFile.scala 71:28]
  reg [31:0] medeleg_data; // @[CsrFile.scala 72:28]
  reg [31:0] mideleg_data; // @[CsrFile.scala 73:28]
  reg [31:0] mepc_data; // @[CsrFile.scala 74:28]
  reg  satp_mode; // @[CsrFile.scala 75:28]
  reg [21:0] satp_ppn; // @[CsrFile.scala 75:28]
  reg [31:0] mtval_data; // @[CsrFile.scala 76:28]
  reg [63:0] mcycle_data; // @[CsrFile.scala 77:28]
  wire [31:0] _T = {mcause_int,mcause_code}; // @[CsrFile.scala 88:49]
  wire [10:0] lo = {2'h0,mstatus_spp,mstatus_mpie,1'h0,mstatus_spie,1'h0,mstatus_mie,1'h0,mstatus_sie,1'h0}; // @[CsrFile.scala 89:50]
  wire [31:0] _T_1 = {13'h0,mstatus_sum,1'h0,2'h0,2'h0,mstatus_mpp,lo}; // @[CsrFile.scala 89:50]
  wire [31:0] _T_2 = {mtvec_base,mtvec_mode}; // @[CsrFile.scala 90:48]
  wire [31:0] _T_3 = {satp_mode,9'h0,satp_ppn}; // @[CsrFile.scala 94:47]
  wire  _T_7 = 12'hf14 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_9 = 12'h342 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_13 = 12'h305 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_15 = 12'h302 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_17 = 12'h303 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_19 = 12'h341 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_21 = 12'h180 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_23 = 12'h343 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_25 = 12'hb00 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_27 = 12'hb80 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_29 = 12'h3a0 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_31 = 12'h3a1 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_33 = 12'h3a2 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_35 = 12'h3a3 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_37 = 12'h3b0 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_39 = 12'h3b1 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_41 = 12'h3b2 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_43 = 12'h3b3 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_45 = 12'h3b4 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_47 = 12'h3b5 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_49 = 12'h3b6 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_51 = 12'h3b7 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_53 = 12'h3b8 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_55 = 12'h3b9 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_57 = 12'h3ba == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_59 = 12'h3bb == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_61 = 12'h3bc == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_63 = 12'h3bd == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_65 = 12'h3be == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_67 = 12'h3bf == io_read_addr; // @[Lookup.scala 31:38]
  wire [31:0] _T_88 = _T_27 ? mcycle_data[63:32] : 32'h0; // @[Lookup.scala 34:39]
  wire [31:0] _T_89 = _T_25 ? mcycle_data[31:0] : _T_88; // @[Lookup.scala 34:39]
  wire [31:0] _T_90 = _T_23 ? mtval_data : _T_89; // @[Lookup.scala 34:39]
  wire [31:0] _T_91 = _T_21 ? _T_3 : _T_90; // @[Lookup.scala 34:39]
  wire [31:0] _T_92 = _T_19 ? mepc_data : _T_91; // @[Lookup.scala 34:39]
  wire [31:0] _T_93 = _T_17 ? mideleg_data : _T_92; // @[Lookup.scala 34:39]
  wire [31:0] _T_94 = _T_15 ? medeleg_data : _T_93; // @[Lookup.scala 34:39]
  wire [31:0] _T_95 = _T_13 ? _T_2 : _T_94; // @[Lookup.scala 34:39]
  wire [31:0] _T_96 = _T_9 ? _T_1 : _T_95; // @[Lookup.scala 34:39]
  wire [31:0] _T_97 = _T_9 ? _T : _T_96; // @[Lookup.scala 34:39]
  wire  readable = _T_7 | (_T_9 | (_T_9 | (_T_13 | (_T_15 | (_T_17 | (_T_19 | (_T_21 | (_T_23 | (_T_25 | (_T_27 | (_T_29
     | (_T_31 | (_T_33 | (_T_35 | (_T_37 | (_T_39 | (_T_41 | (_T_43 | (_T_45 | (_T_47 | (_T_49 | (_T_51 | (_T_53 | (
    _T_55 | (_T_57 | (_T_59 | (_T_61 | (_T_63 | (_T_65 | _T_67))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  writable = _T_7 ? 1'h0 : _T_9 | (_T_9 | (_T_13 | (_T_15 | (_T_17 | (_T_19 | (_T_21 | (_T_23 | (_T_25 | (_T_27 |
    (_T_29 | (_T_31 | (_T_33 | (_T_35 | (_T_37 | (_T_39 | (_T_41 | (_T_43 | (_T_45 | (_T_47 | (_T_49 | (_T_51 | (_T_53
     | (_T_55 | (_T_57 | (_T_59 | (_T_61 | (_T_63 | (_T_65 | _T_67)))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _readValid_T = readable & writable; // @[CsrFile.scala 130:30]
  wire  _readValid_T_6 = 3'h2 == io_read_op ? writable : 3'h1 == io_read_op & readable; // @[Mux.scala 81:58]
  wire  _readValid_T_8 = 3'h3 == io_read_op ? _readValid_T : _readValid_T_6; // @[Mux.scala 81:58]
  wire  _readValid_T_10 = 3'h4 == io_read_op ? _readValid_T : _readValid_T_8; // @[Mux.scala 81:58]
  wire  _csrData_T_1 = 12'hf14 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_3 = 12'h342 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_7 = 12'h305 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_9 = 12'h302 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_11 = 12'h303 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_13 = 12'h341 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_15 = 12'h180 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_17 = 12'h343 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_19 = 12'hb00 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _csrData_T_21 = 12'hb80 == io_write_addr; // @[Lookup.scala 31:38]
  wire [31:0] _csrData_T_82 = _csrData_T_21 ? mcycle_data[63:32] : 32'h0; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_83 = _csrData_T_19 ? mcycle_data[31:0] : _csrData_T_82; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_84 = _csrData_T_17 ? mtval_data : _csrData_T_83; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_85 = _csrData_T_15 ? _T_3 : _csrData_T_84; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_86 = _csrData_T_13 ? mepc_data : _csrData_T_85; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_87 = _csrData_T_11 ? mideleg_data : _csrData_T_86; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_88 = _csrData_T_9 ? medeleg_data : _csrData_T_87; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_89 = _csrData_T_7 ? _T_2 : _csrData_T_88; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_90 = _csrData_T_3 ? _T_1 : _csrData_T_89; // @[Lookup.scala 34:39]
  wire [31:0] _csrData_T_91 = _csrData_T_3 ? _T : _csrData_T_90; // @[Lookup.scala 34:39]
  wire [31:0] csrData = _csrData_T_1 ? 32'h0 : _csrData_T_91; // @[Lookup.scala 34:39]
  wire  writeEn = io_write_op != 3'h0 & io_write_op != 3'h1; // @[CsrFile.scala 140:43]
  wire [31:0] _writeData_T = csrData | io_write_data; // @[CsrFile.scala 144:29]
  wire [31:0] _writeData_T_1 = ~io_write_data; // @[CsrFile.scala 145:31]
  wire [31:0] _writeData_T_2 = csrData & _writeData_T_1; // @[CsrFile.scala 145:29]
  wire [31:0] _writeData_T_4 = 3'h2 == io_write_op ? io_write_data : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _writeData_T_6 = 3'h3 == io_write_op ? io_write_data : _writeData_T_4; // @[Mux.scala 81:58]
  wire [31:0] _writeData_T_8 = 3'h4 == io_write_op ? _writeData_T : _writeData_T_6; // @[Mux.scala 81:58]
  wire [31:0] writeData = 3'h5 == io_write_op ? _writeData_T_2 : _writeData_T_8; // @[Mux.scala 81:58]
  wire [63:0] _mcycle_data_T_1 = mcycle_data + 64'h1; // @[CsrFile.scala 148:32]
  wire [6:0] medeleg_data_lo = {writeData[6],1'h0,writeData[4:2],1'h0,writeData[0]}; // @[Cat.scala 33:92]
  wire [15:0] _medeleg_data_T_6 = {writeData[15],1'h0,writeData[13:12],2'h0,writeData[9:8],1'h0,medeleg_data_lo}; // @[Cat.scala 33:92]
  wire [11:0] _mideleg_data_T_3 = {2'h0,writeData[9],3'h0,writeData[5],3'h0,writeData[1],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] _mepc_data_T_1 = {writeData[31:2],2'h0}; // @[Cat.scala 33:92]
  wire [63:0] _mcycle_data_T_3 = {mcycle_data[63:32],writeData}; // @[Cat.scala 33:92]
  wire [63:0] _mcycle_data_T_5 = {writeData,mcycle_data[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_0 = _csrData_T_21 ? _mcycle_data_T_5 : _mcycle_data_T_1; // @[CsrFile.scala 148:17 151:31 160:43]
  wire [63:0] _GEN_1 = _csrData_T_19 ? _mcycle_data_T_3 : _GEN_0; // @[CsrFile.scala 151:31 159:43]
  wire  _GEN_2 = _csrData_T_15 ? writeData[31] : satp_mode; // @[CsrFile.scala 151:31 CSR.scala 187:11 CsrFile.scala 75:28]
  wire [21:0] _GEN_3 = _csrData_T_15 ? writeData[21:0] : satp_ppn; // @[CsrFile.scala 151:31 CSR.scala 188:11 CsrFile.scala 75:28]
  wire [63:0] _GEN_4 = _csrData_T_15 ? _mcycle_data_T_1 : _GEN_1; // @[CsrFile.scala 148:17 151:31]
  wire [31:0] _GEN_5 = _csrData_T_13 ? _mepc_data_T_1 : mepc_data; // @[CsrFile.scala 151:31 CSR.scala 369:11 CsrFile.scala 74:28]
  wire  _GEN_6 = _csrData_T_13 ? satp_mode : _GEN_2; // @[CsrFile.scala 151:31 75:28]
  wire [21:0] _GEN_7 = _csrData_T_13 ? satp_ppn : _GEN_3; // @[CsrFile.scala 151:31 75:28]
  wire [63:0] _GEN_8 = _csrData_T_13 ? _mcycle_data_T_1 : _GEN_4; // @[CsrFile.scala 148:17 151:31]
  wire [31:0] _GEN_9 = _csrData_T_11 ? {{20'd0}, _mideleg_data_T_3} : mideleg_data; // @[CsrFile.scala 151:31 CSR.scala 271:11 CsrFile.scala 73:28]
  wire [31:0] _GEN_10 = _csrData_T_11 ? mepc_data : _GEN_5; // @[CsrFile.scala 151:31 74:28]
  wire  _GEN_11 = _csrData_T_11 ? satp_mode : _GEN_6; // @[CsrFile.scala 151:31 75:28]
  wire [21:0] _GEN_12 = _csrData_T_11 ? satp_ppn : _GEN_7; // @[CsrFile.scala 151:31 75:28]
  wire [63:0] _GEN_13 = _csrData_T_11 ? _mcycle_data_T_1 : _GEN_8; // @[CsrFile.scala 148:17 151:31]
  wire [31:0] _GEN_14 = _csrData_T_9 ? {{16'd0}, _medeleg_data_T_6} : medeleg_data; // @[CsrFile.scala 151:31 CSR.scala 256:11 CsrFile.scala 72:28]
  wire [31:0] _GEN_15 = _csrData_T_9 ? mideleg_data : _GEN_9; // @[CsrFile.scala 151:31 73:28]
  wire [31:0] _GEN_16 = _csrData_T_9 ? mepc_data : _GEN_10; // @[CsrFile.scala 151:31 74:28]
  wire  _GEN_17 = _csrData_T_9 ? satp_mode : _GEN_11; // @[CsrFile.scala 151:31 75:28]
  wire [21:0] _GEN_18 = _csrData_T_9 ? satp_ppn : _GEN_12; // @[CsrFile.scala 151:31 75:28]
  wire [63:0] _GEN_19 = _csrData_T_9 ? _mcycle_data_T_1 : _GEN_13; // @[CsrFile.scala 148:17 151:31]
  wire [29:0] _GEN_20 = _csrData_T_7 ? writeData[31:2] : mtvec_base; // @[CsrFile.scala 151:31 CSR.scala 345:11 CsrFile.scala 71:28]
  wire [1:0] _GEN_21 = _csrData_T_7 ? {{1'd0}, writeData[0]} : mtvec_mode; // @[CsrFile.scala 151:31 CSR.scala 346:11 CsrFile.scala 71:28]
  wire [31:0] _GEN_22 = _csrData_T_7 ? medeleg_data : _GEN_14; // @[CsrFile.scala 151:31 72:28]
  wire [31:0] _GEN_23 = _csrData_T_7 ? mideleg_data : _GEN_15; // @[CsrFile.scala 151:31 73:28]
  wire [31:0] _GEN_24 = _csrData_T_7 ? mepc_data : _GEN_16; // @[CsrFile.scala 151:31 74:28]
  wire  _GEN_25 = _csrData_T_7 ? satp_mode : _GEN_17; // @[CsrFile.scala 151:31 75:28]
  wire [21:0] _GEN_26 = _csrData_T_7 ? satp_ppn : _GEN_18; // @[CsrFile.scala 151:31 75:28]
  wire [63:0] _GEN_27 = _csrData_T_7 ? _mcycle_data_T_1 : _GEN_19; // @[CsrFile.scala 148:17 151:31]
  wire [31:0] _T_167 = {1'h0,io_except_bits_excCause}; // @[Cat.scala 33:92]
  wire [31:0] _mepc_data_T_3 = {io_except_bits_excPc[31:2],2'h0}; // @[Cat.scala 33:92]
  wire [31:0] csrState_mcycle = mcycle_data[31:0]; // @[CsrFile.scala 179:29]
  wire [31:0] csrState_mcycleh = mcycle_data[63:32]; // @[CsrFile.scala 180:30]
  assign io_read_valid = 3'h5 == io_read_op ? _readValid_T : _readValid_T_10; // @[Mux.scala 81:58]
  assign io_read_data = _T_7 ? 32'h0 : _T_97; // @[Lookup.scala 34:39]
  assign io_mode = 2'h3; // @[CsrFile.scala 171:13]
  assign io_busy = io_write_op != 3'h0 & io_write_op != 3'h1; // @[CsrFile.scala 140:43]
  assign io_mepc = mepc_data; // @[CsrFile.scala 173:13]
  assign io_trapVec = {mtvec_base,mtvec_mode}; // @[CsrFile.scala 174:25]
  assign csrState_0_mcycle = csrState_mcycle;
  assign csrState_0_mcycleh = csrState_mcycleh;
  always @(posedge clock) begin
    if (reset) begin // @[CsrFile.scala 69:28]
      mcause_int <= 1'h0; // @[CsrFile.scala 69:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (_csrData_T_3) begin // @[CsrFile.scala 151:31]
        mcause_int <= writeData[31]; // @[CSR.scala 384:11]
      end
    end else if (io_except_valid) begin // @[CsrFile.scala 162:33]
      mcause_int <= _T_167[31]; // @[CSR.scala 384:11]
    end
    if (reset) begin // @[CsrFile.scala 69:28]
      mcause_code <= 31'h0; // @[CsrFile.scala 69:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (_csrData_T_3) begin // @[CsrFile.scala 151:31]
        mcause_code <= {{27'd0}, writeData[3:0]}; // @[CSR.scala 385:11]
      end
    end else if (io_except_valid) begin // @[CsrFile.scala 162:33]
      mcause_code <= {{27'd0}, _T_167[3:0]}; // @[CSR.scala 385:11]
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_sum <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_sum <= writeData[18]; // @[CSR.scala 222:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_mpp <= 2'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_mpp <= writeData[12:11]; // @[CSR.scala 223:11]
        end
      end
    end else if (io_except_valid) begin // @[CsrFile.scala 162:33]
      mstatus_mpp <= 2'h3; // @[CsrFile.scala 168:22]
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_spp <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_spp <= writeData[8]; // @[CSR.scala 224:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_mpie <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_mpie <= writeData[7]; // @[CSR.scala 225:11]
        end
      end
    end else if (io_except_valid) begin // @[CsrFile.scala 162:33]
      mstatus_mpie <= mstatus_mie; // @[CsrFile.scala 166:22]
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_spie <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_spie <= writeData[5]; // @[CSR.scala 226:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_mie <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_mie <= writeData[3]; // @[CSR.scala 227:11]
        end
      end
    end else if (io_except_valid) begin // @[CsrFile.scala 162:33]
      mstatus_mie <= 1'h0; // @[CsrFile.scala 167:22]
    end
    if (reset) begin // @[CsrFile.scala 70:28]
      mstatus_sie <= 1'h0; // @[CsrFile.scala 70:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
          mstatus_sie <= writeData[1]; // @[CSR.scala 228:11]
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 71:28]
      mtvec_base <= 30'h0; // @[CsrFile.scala 71:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          mtvec_base <= _GEN_20;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 71:28]
      mtvec_mode <= 2'h0; // @[CsrFile.scala 71:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          mtvec_mode <= _GEN_21;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 72:28]
      medeleg_data <= 32'h0; // @[CsrFile.scala 72:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          medeleg_data <= _GEN_22;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 73:28]
      mideleg_data <= 32'h0; // @[CsrFile.scala 73:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          mideleg_data <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 74:28]
      mepc_data <= 32'h0; // @[CsrFile.scala 74:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          mepc_data <= _GEN_24;
        end
      end
    end else if (io_except_valid) begin // @[CsrFile.scala 162:33]
      mepc_data <= _mepc_data_T_3; // @[CSR.scala 369:11]
    end
    if (reset) begin // @[CsrFile.scala 75:28]
      satp_mode <= 1'h0; // @[CsrFile.scala 75:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          satp_mode <= _GEN_25;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 75:28]
      satp_ppn <= 22'h0; // @[CsrFile.scala 75:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (!(_csrData_T_3)) begin // @[CsrFile.scala 151:31]
        if (!(12'h300 == io_write_addr)) begin // @[CsrFile.scala 151:31]
          satp_ppn <= _GEN_26;
        end
      end
    end
    if (reset) begin // @[CsrFile.scala 76:28]
      mtval_data <= 32'h0; // @[CsrFile.scala 76:28]
    end else if (!(writeEn)) begin // @[CsrFile.scala 150:19]
      if (io_except_valid) begin // @[CsrFile.scala 162:33]
        mtval_data <= io_except_bits_excValue; // @[CSR.scala 17:10]
      end
    end
    if (reset) begin // @[CsrFile.scala 77:28]
      mcycle_data <= 64'h0; // @[CsrFile.scala 77:28]
    end else if (writeEn) begin // @[CsrFile.scala 150:19]
      if (_csrData_T_3) begin // @[CsrFile.scala 151:31]
        mcycle_data <= _mcycle_data_T_1; // @[CsrFile.scala 148:17]
      end else if (12'h300 == io_write_addr) begin // @[CsrFile.scala 151:31]
        mcycle_data <= _mcycle_data_T_1; // @[CsrFile.scala 148:17]
      end else begin
        mcycle_data <= _GEN_27;
      end
    end else begin
      mcycle_data <= _mcycle_data_T_1; // @[CsrFile.scala 148:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mcause_int = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mcause_code = _RAND_1[30:0];
  _RAND_2 = {1{`RANDOM}};
  mstatus_sum = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  mstatus_mpp = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  mstatus_spp = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  mstatus_mpie = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  mstatus_spie = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  mstatus_mie = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mstatus_sie = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  mtvec_base = _RAND_9[29:0];
  _RAND_10 = {1{`RANDOM}};
  mtvec_mode = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  medeleg_data = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mideleg_data = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mepc_data = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  satp_mode = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  satp_ppn = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  mtval_data = _RAND_16[31:0];
  _RAND_17 = {2{`RANDOM}};
  mcycle_data = _RAND_17[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBusArbiter(
  input        clock,
  input        reset,
  input        io_reqs_1,
  output [1:0] io_grantOH
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] owner; // @[Bus.scala 162:24]
  wire [3:0] _io_grantOH_T = 4'h1 << owner; // @[OneHot.scala 57:35]
  assign io_grantOH = _io_grantOH_T[1:0]; // @[Bus.scala 190:16]
  always @(posedge clock) begin
    if (reset) begin // @[Bus.scala 162:24]
      owner <= 2'h0; // @[Bus.scala 162:24]
    end else if (io_reqs_1) begin // @[Mux.scala 27:73]
      owner <= 2'h1;
    end else begin
      owner <= 2'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  owner = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBusMux(
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [31:0]  io_in_0_bits_address,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [2:0]   io_in_1_bits_opcode,
  input  [31:0]  io_in_1_bits_address,
  input  [127:0] io_in_1_bits_data,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_opcode,
  output [127:0] io_out_bits_size,
  output         io_out_bits_source,
  output [31:0]  io_out_bits_address,
  output [127:0] io_out_bits_data,
  input          io_choseOH_0,
  input          io_choseOH_1
);
  wire [31:0] _io_out_bits_T_9 = io_choseOH_0 ? io_in_0_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_bits_T_10 = io_choseOH_1 ? io_in_1_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [127:0] _io_out_bits_T_15 = io_choseOH_0 ? 128'h20 : 128'h0; // @[Mux.scala 27:73]
  wire [127:0] _io_out_bits_T_16 = io_choseOH_1 ? 128'h10 : 128'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_21 = io_choseOH_0 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_22 = io_choseOH_1 ? io_in_1_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  assign io_in_0_ready = io_out_ready & io_choseOH_0; // @[Bus.scala 132:80]
  assign io_in_1_ready = io_out_ready & io_choseOH_1; // @[Bus.scala 132:80]
  assign io_out_valid = io_choseOH_0 & io_in_0_valid | io_choseOH_1 & io_in_1_valid; // @[Mux.scala 27:73]
  assign io_out_bits_opcode = _io_out_bits_T_21 | _io_out_bits_T_22; // @[Mux.scala 27:73]
  assign io_out_bits_size = _io_out_bits_T_15 | _io_out_bits_T_16; // @[Mux.scala 27:73]
  assign io_out_bits_source = io_choseOH_1; // @[Mux.scala 27:73]
  assign io_out_bits_address = _io_out_bits_T_9 | _io_out_bits_T_10; // @[Mux.scala 27:73]
  assign io_out_bits_data = io_choseOH_1 ? io_in_1_bits_data : 128'h0; // @[Mux.scala 27:73]
endmodule
module Queue(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [2:0]   io_enq_bits_opcode,
  input  [127:0] io_enq_bits_size,
  input          io_enq_bits_source,
  input  [31:0]  io_enq_bits_address,
  input  [127:0] io_enq_bits_data,
  input          io_deq_ready,
  output         io_deq_valid,
  output [2:0]   io_deq_bits_opcode,
  output [127:0] io_deq_bits_size,
  output         io_deq_bits_source,
  output [31:0]  io_deq_bits_address,
  output [127:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_opcode_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 273:95]
  reg [127:0] ram_size [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [127:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [127:0] ram_size_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_source [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg [31:0] ram_address [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_address_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 273:95]
  reg [127:0] ram_data [0:7]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [2:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [127:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [127:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire  _GEN_19 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_19 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = enq_ptr_value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_19 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_opcode = empty ? io_enq_bits_opcode : ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_source = empty ? io_enq_bits_source : ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_address = empty ? io_enq_bits_address : ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[127:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_address[initvar] = _RAND_3[31:0];
  _RAND_4 = {4{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_data[initvar] = _RAND_4[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enq_ptr_value = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  deq_ptr_value = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLAddrDecode(
  input  [31:0] io_addr,
  output        io_choseOH_0,
  output        io_choseOH_1
);
  wire  valid = io_addr < 32'h10000000; // @[Bus.scala 201:42]
  wire  valid_1 = io_addr >= 32'h10000000 & io_addr < 32'h20000000; // @[Bus.scala 201:31]
  wire  _GEN_2 = valid_1 ? 1'h0 : 1'h1; // @[Bus.scala 211:68 212:20 214:20]
  assign io_choseOH_0 = valid | _GEN_2; // @[Bus.scala 209:62 210:20]
  assign io_choseOH_1 = valid ? 1'h0 : valid_1; // @[Bus.scala 209:62 210:20]
endmodule
module TLBusMux_1(
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [2:0]   io_in_0_bits_opcode,
  input  [127:0] io_in_0_bits_data,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_opcode,
  output [127:0] io_out_bits_data,
  input          io_choseOH_0
);
  assign io_in_0_ready = io_out_ready & io_choseOH_0; // @[Bus.scala 132:80]
  assign io_out_valid = io_choseOH_0 & io_in_0_valid; // @[Mux.scala 27:73]
  assign io_out_bits_opcode = io_choseOH_0 ? io_in_0_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  assign io_out_bits_data = io_choseOH_0 ? io_in_0_bits_data : 128'h0; // @[Mux.scala 27:73]
endmodule
module TLXbar(
  input          clock,
  input          reset,
  output         io_masterFace_in_0_ready,
  input          io_masterFace_in_0_valid,
  input  [31:0]  io_masterFace_in_0_bits_address,
  output         io_masterFace_in_1_ready,
  input          io_masterFace_in_1_valid,
  input  [2:0]   io_masterFace_in_1_bits_opcode,
  input  [31:0]  io_masterFace_in_1_bits_address,
  input  [127:0] io_masterFace_in_1_bits_data,
  output         io_masterFace_out_0_valid,
  output [2:0]   io_masterFace_out_0_bits_opcode,
  output [127:0] io_masterFace_out_0_bits_data,
  output         io_masterFace_out_1_valid,
  output [2:0]   io_masterFace_out_1_bits_opcode,
  output [127:0] io_masterFace_out_1_bits_data,
  input          io_slaveFace_in_0_ready,
  output         io_slaveFace_in_0_valid,
  output [2:0]   io_slaveFace_in_0_bits_opcode,
  output [127:0] io_slaveFace_in_0_bits_size,
  output [31:0]  io_slaveFace_in_0_bits_address,
  output [127:0] io_slaveFace_in_0_bits_data,
  output         io_slaveFace_out_0_ready,
  input          io_slaveFace_out_0_valid,
  input  [2:0]   io_slaveFace_out_0_bits_opcode,
  input  [127:0] io_slaveFace_out_0_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  reqArb_clock; // @[Bus.scala 233:24]
  wire  reqArb_reset; // @[Bus.scala 233:24]
  wire  reqArb_io_reqs_1; // @[Bus.scala 233:24]
  wire [1:0] reqArb_io_grantOH; // @[Bus.scala 233:24]
  wire  reqMux_io_in_0_ready; // @[Bus.scala 236:24]
  wire  reqMux_io_in_0_valid; // @[Bus.scala 236:24]
  wire [31:0] reqMux_io_in_0_bits_address; // @[Bus.scala 236:24]
  wire  reqMux_io_in_1_ready; // @[Bus.scala 236:24]
  wire  reqMux_io_in_1_valid; // @[Bus.scala 236:24]
  wire [2:0] reqMux_io_in_1_bits_opcode; // @[Bus.scala 236:24]
  wire [31:0] reqMux_io_in_1_bits_address; // @[Bus.scala 236:24]
  wire [127:0] reqMux_io_in_1_bits_data; // @[Bus.scala 236:24]
  wire  reqMux_io_out_ready; // @[Bus.scala 236:24]
  wire  reqMux_io_out_valid; // @[Bus.scala 236:24]
  wire [2:0] reqMux_io_out_bits_opcode; // @[Bus.scala 236:24]
  wire [127:0] reqMux_io_out_bits_size; // @[Bus.scala 236:24]
  wire  reqMux_io_out_bits_source; // @[Bus.scala 236:24]
  wire [31:0] reqMux_io_out_bits_address; // @[Bus.scala 236:24]
  wire [127:0] reqMux_io_out_bits_data; // @[Bus.scala 236:24]
  wire  reqMux_io_choseOH_0; // @[Bus.scala 236:24]
  wire  reqMux_io_choseOH_1; // @[Bus.scala 236:24]
  wire  buf__clock; // @[Bus.scala 242:21]
  wire  buf__reset; // @[Bus.scala 242:21]
  wire  buf__io_enq_ready; // @[Bus.scala 242:21]
  wire  buf__io_enq_valid; // @[Bus.scala 242:21]
  wire [2:0] buf__io_enq_bits_opcode; // @[Bus.scala 242:21]
  wire [127:0] buf__io_enq_bits_size; // @[Bus.scala 242:21]
  wire  buf__io_enq_bits_source; // @[Bus.scala 242:21]
  wire [31:0] buf__io_enq_bits_address; // @[Bus.scala 242:21]
  wire [127:0] buf__io_enq_bits_data; // @[Bus.scala 242:21]
  wire  buf__io_deq_ready; // @[Bus.scala 242:21]
  wire  buf__io_deq_valid; // @[Bus.scala 242:21]
  wire [2:0] buf__io_deq_bits_opcode; // @[Bus.scala 242:21]
  wire [127:0] buf__io_deq_bits_size; // @[Bus.scala 242:21]
  wire  buf__io_deq_bits_source; // @[Bus.scala 242:21]
  wire [31:0] buf__io_deq_bits_address; // @[Bus.scala 242:21]
  wire [127:0] buf__io_deq_bits_data; // @[Bus.scala 242:21]
  wire [31:0] addrDec_io_addr; // @[Bus.scala 265:25]
  wire  addrDec_io_choseOH_0; // @[Bus.scala 265:25]
  wire  addrDec_io_choseOH_1; // @[Bus.scala 265:25]
  wire  slaveMux_io_in_0_ready; // @[Bus.scala 310:26]
  wire  slaveMux_io_in_0_valid; // @[Bus.scala 310:26]
  wire [2:0] slaveMux_io_in_0_bits_opcode; // @[Bus.scala 310:26]
  wire [127:0] slaveMux_io_in_0_bits_data; // @[Bus.scala 310:26]
  wire  slaveMux_io_out_ready; // @[Bus.scala 310:26]
  wire  slaveMux_io_out_valid; // @[Bus.scala 310:26]
  wire [2:0] slaveMux_io_out_bits_opcode; // @[Bus.scala 310:26]
  wire [127:0] slaveMux_io_out_bits_data; // @[Bus.scala 310:26]
  wire  slaveMux_io_choseOH_0; // @[Bus.scala 310:26]
  wire [1:0] _WIRE_1 = reqArb_io_grantOH; // @[Bus.scala 238:{52,52}]
  reg  s1_full; // @[Bus.scala 249:26]
  wire  s1_latch = buf__io_deq_ready & buf__io_deq_valid; // @[Decoupled.scala 51:35]
  reg [2:0] s1_req_opcode; // @[Reg.scala 19:16]
  reg [127:0] s1_req_size; // @[Reg.scala 19:16]
  reg  s1_req_source; // @[Reg.scala 19:16]
  reg [31:0] s1_req_address; // @[Reg.scala 19:16]
  reg [127:0] s1_req_data; // @[Reg.scala 19:16]
  wire [123:0] s1_beatSize = s1_req_size[127:4]; // @[Bus.scala 255:35]
  reg [4:0] s1_beatCounter_value; // @[Counter.scala 61:40]
  wire [123:0] _s1_lastBeat_T_1 = s1_beatSize - 124'h1; // @[Bus.scala 278:60]
  wire [123:0] _GEN_27 = {{119'd0}, s1_beatCounter_value}; // @[Bus.scala 278:44]
  wire  s1_lastBeat = _GEN_27 == _s1_lastBeat_T_1; // @[Bus.scala 278:44]
  wire  _s1_putMultiBeat_T = ~s1_lastBeat; // @[Bus.scala 287:25]
  wire  _s1_putMultiBeat_T_1 = s1_req_opcode == 3'h2; // @[Bus.scala 287:55]
  wire  s1_putMultiBeat = ~s1_lastBeat & s1_req_opcode == 3'h2; // @[Bus.scala 287:38]
  reg  s2_full; // @[Bus.scala 297:26]
  reg [2:0] s2_opcode; // @[Reg.scala 19:16]
  wire [1:0] s2_masterRecvVec = {io_masterFace_out_1_valid,io_masterFace_out_0_valid}; // @[Cat.scala 33:92]
  reg [1:0] s2_chosenMasterOH; // @[Reg.scala 19:16]
  wire [1:0] _s2_masterRecv_T = s2_masterRecvVec & s2_chosenMasterOH; // @[Bus.scala 322:43]
  wire  s2_masterRecv = |_s2_masterRecv_T; // @[Bus.scala 322:64]
  reg  s2_masterRecvHold_holdReg; // @[Reg.scala 19:16]
  wire  s2_masterRecvHold = s2_masterRecv ? s2_masterRecv : s2_masterRecvHold_holdReg; // @[util.scala 26:12]
  reg [4:0] s2_beatCounter_value; // @[Counter.scala 61:40]
  reg [123:0] s2_beatSize; // @[Reg.scala 19:16]
  wire [123:0] _s2_lastBeat_T_1 = s2_beatSize - 124'h1; // @[Bus.scala 324:60]
  wire [123:0] _GEN_28 = {{119'd0}, s2_beatCounter_value}; // @[Bus.scala 324:44]
  wire  s2_lastBeat = _GEN_28 == _s2_lastBeat_T_1; // @[Bus.scala 324:44]
  wire  s2_getAllBeat = s2_opcode == 3'h4 & s2_masterRecvHold & s2_lastBeat; // @[Bus.scala 332:61]
  wire  s2_fire = s2_opcode == 3'h2 & s2_masterRecvHold | s2_getAllBeat; // @[Bus.scala 333:65]
  wire  s2_ready = ~s2_full | s2_fire; // @[Bus.scala 306:26]
  wire  _s1_slaveRecVec_T = io_slaveFace_in_0_ready & io_slaveFace_in_0_valid; // @[Decoupled.scala 51:35]
  wire [1:0] s1_slaveRecVec = {1'h0,_s1_slaveRecVec_T}; // @[Cat.scala 33:92]
  wire [1:0] _s1_slaveRecv_T = {addrDec_io_choseOH_1,addrDec_io_choseOH_0}; // @[Bus.scala 276:59]
  wire [1:0] _s1_slaveRecv_T_1 = s1_slaveRecVec & _s1_slaveRecv_T; // @[Bus.scala 276:40]
  wire  s1_slaveRecv = |_s1_slaveRecv_T_1; // @[Bus.scala 276:67]
  reg  s1_slaveRecvHold_holdReg; // @[Reg.scala 19:16]
  wire  s1_slaveRecvHold = s1_slaveRecv ? s1_slaveRecv : s1_slaveRecvHold_holdReg; // @[util.scala 26:12]
  wire  s1_putAllBeat = s1_lastBeat & _s1_putMultiBeat_T_1; // @[Bus.scala 289:34]
  wire  s1_valid = s1_slaveRecvHold & (s1_putAllBeat | s1_req_opcode == 3'h4); // @[Bus.scala 290:34]
  wire  s1_fire = s2_ready & s1_valid; // @[Bus.scala 292:25]
  wire  _GEN_8 = s1_full & s1_fire ? 1'h0 : s1_full; // @[Bus.scala 249:26 263:{35,45}]
  wire  _GEN_9 = s1_latch | _GEN_8; // @[Bus.scala 262:{20,30}]
  wire [4:0] _value_T_1 = s1_beatCounter_value + 5'h1; // @[Counter.scala 77:24]
  reg  s2_chosenSlaveOH_0; // @[Reg.scala 19:16]
  wire [1:0] _s2_chosenMasterOH_T = 2'h1 << s1_req_source; // @[OneHot.scala 57:35]
  wire  _GEN_19 = s2_full & s2_fire ? 1'h0 : s2_full; // @[Bus.scala 297:26 308:{35,45}]
  wire  _GEN_20 = s1_fire | _GEN_19; // @[Bus.scala 307:{20,30}]
  wire [4:0] _value_T_3 = s2_beatCounter_value + 5'h1; // @[Counter.scala 77:24]
  reg  idle; // @[Bus.scala 337:23]
  wire  _GEN_25 = s2_fire | idle; // @[Bus.scala 341:26 342:14 337:23]
  wire  _GEN_26 = s1_latch | s1_fire ? 1'h0 : _GEN_25; // @[Bus.scala 339:32 340:14]
  TLBusArbiter reqArb ( // @[Bus.scala 233:24]
    .clock(reqArb_clock),
    .reset(reqArb_reset),
    .io_reqs_1(reqArb_io_reqs_1),
    .io_grantOH(reqArb_io_grantOH)
  );
  TLBusMux reqMux ( // @[Bus.scala 236:24]
    .io_in_0_ready(reqMux_io_in_0_ready),
    .io_in_0_valid(reqMux_io_in_0_valid),
    .io_in_0_bits_address(reqMux_io_in_0_bits_address),
    .io_in_1_ready(reqMux_io_in_1_ready),
    .io_in_1_valid(reqMux_io_in_1_valid),
    .io_in_1_bits_opcode(reqMux_io_in_1_bits_opcode),
    .io_in_1_bits_address(reqMux_io_in_1_bits_address),
    .io_in_1_bits_data(reqMux_io_in_1_bits_data),
    .io_out_ready(reqMux_io_out_ready),
    .io_out_valid(reqMux_io_out_valid),
    .io_out_bits_opcode(reqMux_io_out_bits_opcode),
    .io_out_bits_size(reqMux_io_out_bits_size),
    .io_out_bits_source(reqMux_io_out_bits_source),
    .io_out_bits_address(reqMux_io_out_bits_address),
    .io_out_bits_data(reqMux_io_out_bits_data),
    .io_choseOH_0(reqMux_io_choseOH_0),
    .io_choseOH_1(reqMux_io_choseOH_1)
  );
  Queue buf_ ( // @[Bus.scala 242:21]
    .clock(buf__clock),
    .reset(buf__reset),
    .io_enq_ready(buf__io_enq_ready),
    .io_enq_valid(buf__io_enq_valid),
    .io_enq_bits_opcode(buf__io_enq_bits_opcode),
    .io_enq_bits_size(buf__io_enq_bits_size),
    .io_enq_bits_source(buf__io_enq_bits_source),
    .io_enq_bits_address(buf__io_enq_bits_address),
    .io_enq_bits_data(buf__io_enq_bits_data),
    .io_deq_ready(buf__io_deq_ready),
    .io_deq_valid(buf__io_deq_valid),
    .io_deq_bits_opcode(buf__io_deq_bits_opcode),
    .io_deq_bits_size(buf__io_deq_bits_size),
    .io_deq_bits_source(buf__io_deq_bits_source),
    .io_deq_bits_address(buf__io_deq_bits_address),
    .io_deq_bits_data(buf__io_deq_bits_data)
  );
  TLAddrDecode addrDec ( // @[Bus.scala 265:25]
    .io_addr(addrDec_io_addr),
    .io_choseOH_0(addrDec_io_choseOH_0),
    .io_choseOH_1(addrDec_io_choseOH_1)
  );
  TLBusMux_1 slaveMux ( // @[Bus.scala 310:26]
    .io_in_0_ready(slaveMux_io_in_0_ready),
    .io_in_0_valid(slaveMux_io_in_0_valid),
    .io_in_0_bits_opcode(slaveMux_io_in_0_bits_opcode),
    .io_in_0_bits_data(slaveMux_io_in_0_bits_data),
    .io_out_ready(slaveMux_io_out_ready),
    .io_out_valid(slaveMux_io_out_valid),
    .io_out_bits_opcode(slaveMux_io_out_bits_opcode),
    .io_out_bits_data(slaveMux_io_out_bits_data),
    .io_choseOH_0(slaveMux_io_choseOH_0)
  );
  assign io_masterFace_in_0_ready = reqMux_io_in_0_ready; // @[Bus.scala 237:58]
  assign io_masterFace_in_1_ready = reqMux_io_in_1_ready; // @[Bus.scala 237:58]
  assign io_masterFace_out_0_valid = slaveMux_io_out_valid & s2_chosenMasterOH[0]; // @[Bus.scala 316:43]
  assign io_masterFace_out_0_bits_opcode = slaveMux_io_out_bits_opcode; // @[Bus.scala 315:17]
  assign io_masterFace_out_0_bits_data = slaveMux_io_out_bits_data; // @[Bus.scala 315:17]
  assign io_masterFace_out_1_valid = slaveMux_io_out_valid & s2_chosenMasterOH[1]; // @[Bus.scala 316:43]
  assign io_masterFace_out_1_bits_opcode = slaveMux_io_out_bits_opcode; // @[Bus.scala 315:17]
  assign io_masterFace_out_1_bits_data = slaveMux_io_out_bits_data; // @[Bus.scala 315:17]
  assign io_slaveFace_in_0_valid = addrDec_io_choseOH_0 & s1_full; // @[Bus.scala 271:41]
  assign io_slaveFace_in_0_bits_opcode = s1_req_opcode; // @[Bus.scala 270:18]
  assign io_slaveFace_in_0_bits_size = s1_req_size; // @[Bus.scala 270:18]
  assign io_slaveFace_in_0_bits_address = s1_req_address; // @[Bus.scala 270:18]
  assign io_slaveFace_in_0_bits_data = s1_req_data; // @[Bus.scala 270:18]
  assign io_slaveFace_out_0_ready = slaveMux_io_in_0_ready; // @[Bus.scala 311:20]
  assign reqArb_clock = clock;
  assign reqArb_reset = reset;
  assign reqArb_io_reqs_1 = io_masterFace_in_1_valid; // @[Bus.scala 234:58]
  assign reqMux_io_in_0_valid = io_masterFace_in_0_valid; // @[Bus.scala 237:58]
  assign reqMux_io_in_0_bits_address = io_masterFace_in_0_bits_address; // @[Bus.scala 237:58]
  assign reqMux_io_in_1_valid = io_masterFace_in_1_valid; // @[Bus.scala 237:58]
  assign reqMux_io_in_1_bits_opcode = io_masterFace_in_1_bits_opcode; // @[Bus.scala 237:58]
  assign reqMux_io_in_1_bits_address = io_masterFace_in_1_bits_address; // @[Bus.scala 237:58]
  assign reqMux_io_in_1_bits_data = io_masterFace_in_1_bits_data; // @[Bus.scala 237:58]
  assign reqMux_io_out_ready = buf__io_enq_ready; // @[Bus.scala 243:16]
  assign reqMux_io_choseOH_0 = _WIRE_1[0]; // @[Bus.scala 238:52]
  assign reqMux_io_choseOH_1 = _WIRE_1[1]; // @[Bus.scala 238:52]
  assign buf__clock = clock;
  assign buf__reset = reset;
  assign buf__io_enq_valid = reqMux_io_out_valid; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_opcode = reqMux_io_out_bits_opcode; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_size = reqMux_io_out_bits_size; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_source = reqMux_io_out_bits_source; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_address = reqMux_io_out_bits_address; // @[Bus.scala 243:16]
  assign buf__io_enq_bits_data = reqMux_io_out_bits_data; // @[Bus.scala 243:16]
  assign buf__io_deq_ready = ~s1_full | s1_putMultiBeat | s1_fire; // @[Bus.scala 261:45]
  assign addrDec_io_addr = s1_req_address; // @[Bus.scala 267:21]
  assign slaveMux_io_in_0_valid = io_slaveFace_out_0_valid; // @[Bus.scala 311:20]
  assign slaveMux_io_in_0_bits_opcode = io_slaveFace_out_0_bits_opcode; // @[Bus.scala 311:20]
  assign slaveMux_io_in_0_bits_data = io_slaveFace_out_0_bits_data; // @[Bus.scala 311:20]
  assign slaveMux_io_out_ready = s2_chosenMasterOH[0] | s2_chosenMasterOH[1]; // @[Mux.scala 27:73]
  assign slaveMux_io_choseOH_0 = s2_chosenSlaveOH_0; // @[Bus.scala 312:25]
  always @(posedge clock) begin
    if (reset) begin // @[Bus.scala 249:26]
      s1_full <= 1'h0; // @[Bus.scala 249:26]
    end else begin
      s1_full <= _GEN_9;
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_opcode <= buf__io_deq_bits_opcode; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_size <= buf__io_deq_bits_size; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_source <= buf__io_deq_bits_source; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_address <= buf__io_deq_bits_address; // @[Reg.scala 20:22]
    end
    if (s1_latch) begin // @[Reg.scala 20:18]
      s1_req_data <= buf__io_deq_bits_data; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Counter.scala 61:40]
      s1_beatCounter_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (s1_fire) begin // @[Bus.scala 282:19]
      s1_beatCounter_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (s1_slaveRecv & _s1_putMultiBeat_T) begin // @[Bus.scala 279:40]
      s1_beatCounter_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Bus.scala 297:26]
      s2_full <= 1'h0; // @[Bus.scala 297:26]
    end else begin
      s2_full <= _GEN_20;
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_opcode <= s1_req_opcode; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_chosenMasterOH <= _s2_chosenMasterOH_T; // @[Reg.scala 20:22]
    end
    if (s2_fire) begin // @[util.scala 25:21]
      s2_masterRecvHold_holdReg <= 1'h0; // @[util.scala 25:31]
    end else if (s2_masterRecv) begin // @[util.scala 26:12]
      s2_masterRecvHold_holdReg <= s2_masterRecv;
    end
    if (reset) begin // @[Counter.scala 61:40]
      s2_beatCounter_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (s2_fire) begin // @[Bus.scala 328:19]
      s2_beatCounter_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (s2_masterRecv & ~s2_lastBeat) begin // @[Bus.scala 325:41]
      s2_beatCounter_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_beatSize <= s1_beatSize; // @[Reg.scala 20:22]
    end
    if (s1_fire) begin // @[util.scala 25:21]
      s1_slaveRecvHold_holdReg <= 1'h0; // @[util.scala 25:31]
    end else if (s1_slaveRecv) begin // @[util.scala 26:12]
      s1_slaveRecvHold_holdReg <= s1_slaveRecv;
    end
    if (s1_fire) begin // @[Reg.scala 20:18]
      s2_chosenSlaveOH_0 <= addrDec_io_choseOH_0; // @[Reg.scala 20:22]
    end
    idle <= reset | _GEN_26; // @[Bus.scala 337:{23,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s1_req_opcode = _RAND_1[2:0];
  _RAND_2 = {4{`RANDOM}};
  s1_req_size = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  s1_req_source = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s1_req_address = _RAND_4[31:0];
  _RAND_5 = {4{`RANDOM}};
  s1_req_data = _RAND_5[127:0];
  _RAND_6 = {1{`RANDOM}};
  s1_beatCounter_value = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  s2_full = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s2_opcode = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  s2_chosenMasterOH = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  s2_masterRecvHold_holdReg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  s2_beatCounter_value = _RAND_11[4:0];
  _RAND_12 = {4{`RANDOM}};
  s2_beatSize = _RAND_12[123:0];
  _RAND_13 = {1{`RANDOM}};
  s1_slaveRecvHold_holdReg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  s2_chosenSlaveOH_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  idle = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SingleROM(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [2:0]   io_req_bits_opcode,
  input  [127:0] io_req_bits_size,
  input  [31:0]  io_req_bits_address,
  input  [127:0] io_req_bits_data,
  input          io_resp_ready,
  output         io_resp_valid,
  output [2:0]   io_resp_bits_opcode,
  output [127:0] io_resp_bits_size,
  output [127:0] io_resp_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] mem [0:131071]; // @[SingleROM.scala 14:26]
  wire  mem_rdata_en; // @[SingleROM.scala 14:26]
  wire [16:0] mem_rdata_addr; // @[SingleROM.scala 14:26]
  wire [127:0] mem_rdata_data; // @[SingleROM.scala 14:26]
  wire [127:0] mem_MPORT_data; // @[SingleROM.scala 14:26]
  wire [16:0] mem_MPORT_addr; // @[SingleROM.scala 14:26]
  wire  mem_MPORT_mask; // @[SingleROM.scala 14:26]
  wire  mem_MPORT_en; // @[SingleROM.scala 14:26]
  reg  mem_rdata_en_pipe_0;
  reg [16:0] mem_rdata_addr_pipe_0;
  wire  _reqReg_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  reg [2:0] reqReg_opcode; // @[Reg.scala 19:16]
  reg [127:0] reqReg_size; // @[Reg.scala 19:16]
  reg [31:0] reqReg_address; // @[Reg.scala 19:16]
  reg [127:0] reqReg_data; // @[Reg.scala 19:16]
  wire [2:0] _GEN_0 = _reqReg_T ? io_req_bits_opcode : reqReg_opcode; // @[Reg.scala 19:16 20:{18,22}]
  wire [31:0] _GEN_4 = _reqReg_T ? io_req_bits_address : reqReg_address; // @[Reg.scala 19:16 20:{18,22}]
  reg  busy; // @[SingleROM.scala 19:23]
  reg [4:0] reqLastBeat_count_value; // @[Counter.scala 61:40]
  wire [123:0] reqLastBeat_beatNum = io_req_bits_size[127:4]; // @[Bus.scala 85:41]
  wire [123:0] _reqLastBeat_lastBeat_T_1 = reqLastBeat_beatNum - 124'h1; // @[Bus.scala 86:52]
  wire [123:0] _GEN_25 = {{119'd0}, reqLastBeat_count_value}; // @[Bus.scala 86:40]
  wire  reqLastBeat_lastBeat = _GEN_25 == _reqLastBeat_lastBeat_T_1; // @[Bus.scala 86:40]
  wire  reqLastBeat_fireLastBeat = _reqReg_T & reqLastBeat_lastBeat; // @[Bus.scala 87:38]
  wire [4:0] _reqLastBeat_value_T_1 = reqLastBeat_count_value + 5'h1; // @[Counter.scala 77:24]
  reg [4:0] respLastBeat_count_value; // @[Counter.scala 61:40]
  wire [123:0] respLastBeat_beatNum = io_resp_bits_size[127:4]; // @[Bus.scala 96:42]
  wire [123:0] _respLastBeat_lastBeat_T_1 = respLastBeat_beatNum - 124'h1; // @[Bus.scala 97:52]
  wire [123:0] _GEN_26 = {{119'd0}, respLastBeat_count_value}; // @[Bus.scala 97:40]
  wire  respLastBeat_lastBeat = _GEN_26 == _respLastBeat_lastBeat_T_1; // @[Bus.scala 97:40]
  wire  _respLastBeat_fireLastBeat_T = io_resp_ready & io_resp_valid; // @[Decoupled.scala 51:35]
  wire  respLastBeat_fireLastBeat = _respLastBeat_fireLastBeat_T & respLastBeat_lastBeat; // @[Bus.scala 98:39]
  wire [4:0] _respLastBeat_value_T_1 = respLastBeat_count_value + 5'h1; // @[Counter.scala 77:24]
  wire  _getFire_T_1 = _GEN_0 == 3'h4; // @[SingleROM.scala 27:45]
  wire  getFire = _reqReg_T & _GEN_0 == 3'h4; // @[SingleROM.scala 27:31]
  wire  _putFire_T_2 = _GEN_0 == 3'h2; // @[SingleROM.scala 28:60]
  wire  putFire = _reqReg_T & reqLastBeat_fireLastBeat & _GEN_0 == 3'h2; // @[SingleROM.scala 28:46]
  wire  reqLatch = getFire | putFire; // @[SingleROM.scala 29:28]
  wire  _finish_T_2 = reqReg_opcode == 3'h4; // @[SingleROM.scala 58:86]
  wire  finish = _respLastBeat_fireLastBeat_T & (reqReg_opcode == 3'h2 | reqReg_opcode == 3'h4 &
    respLastBeat_fireLastBeat); // @[SingleROM.scala 58:28]
  wire  _GEN_12 = busy & finish ? 1'h0 : busy; // @[SingleROM.scala 19:23 31:{31,38}]
  wire  _GEN_13 = reqLatch | _GEN_12; // @[SingleROM.scala 30:{20,27}]
  wire  ren = _getFire_T_1 & (_reqReg_T | _respLastBeat_fireLastBeat_T); // @[SingleROM.scala 33:41]
  wire  wen = _reqReg_T & _putFire_T_2; // @[SingleROM.scala 34:27]
  reg [4:0] beatCount_count_value; // @[Counter.scala 61:40]
  wire [123:0] _GEN_27 = {{119'd0}, beatCount_count_value}; // @[Bus.scala 97:40]
  wire  beatCount_lastBeat = _GEN_27 == _respLastBeat_lastBeat_T_1; // @[Bus.scala 97:40]
  wire  beatCount_fireLastBeat = _respLastBeat_fireLastBeat_T & beatCount_lastBeat; // @[Bus.scala 98:39]
  wire [4:0] _beatCount_value_T_1 = beatCount_count_value + 5'h1; // @[Counter.scala 77:24]
  wire [4:0] beatCount = _reqReg_T ? 5'h0 : _beatCount_value_T_1; // @[SingleROM.scala 38:24]
  wire [8:0] addrOff = {beatCount, 4'h0}; // @[SingleROM.scala 39:29]
  wire [31:0] _GEN_28 = {{23'd0}, addrOff}; // @[SingleROM.scala 40:31]
  wire [31:0] _rdAddr_T_1 = _GEN_4 + _GEN_28; // @[SingleROM.scala 40:31]
  wire [27:0] rdAddr = _rdAddr_T_1[31:4]; // @[SingleROM.scala 40:42]
  wire [27:0] wrAddr = _GEN_4[31:4]; // @[SingleROM.scala 45:30]
  assign mem_rdata_en = mem_rdata_en_pipe_0;
  assign mem_rdata_addr = mem_rdata_addr_pipe_0;
  assign mem_rdata_data = mem[mem_rdata_addr]; // @[SingleROM.scala 14:26]
  assign mem_MPORT_data = _reqReg_T ? io_req_bits_data : reqReg_data;
  assign mem_MPORT_addr = wrAddr[16:0];
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = wen;
  assign io_req_ready = ~busy; // @[SingleROM.scala 22:21]
  assign io_resp_valid = busy; // @[SingleROM.scala 51:19]
  assign io_resp_bits_opcode = {{2'd0}, _finish_T_2}; // @[SingleROM.scala 55:25]
  assign io_resp_bits_size = reqReg_size; // @[SingleROM.scala 53:23]
  assign io_resp_bits_data = mem_rdata_data; // @[SingleROM.scala 54:23]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SingleROM.scala 14:26]
    end
    mem_rdata_en_pipe_0 <= ren;
    if (ren) begin
      mem_rdata_addr_pipe_0 <= rdAddr[16:0];
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_opcode <= io_req_bits_opcode; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_size <= io_req_bits_size; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_address <= io_req_bits_address; // @[Reg.scala 20:22]
    end
    if (_reqReg_T) begin // @[Reg.scala 20:18]
      reqReg_data <= io_req_bits_data; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[SingleROM.scala 19:23]
      busy <= 1'h0; // @[SingleROM.scala 19:23]
    end else begin
      busy <= _GEN_13;
    end
    if (reset) begin // @[Counter.scala 61:40]
      reqLastBeat_count_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (reqLastBeat_fireLastBeat | _reqReg_T & io_req_bits_opcode == 3'h4) begin // @[Bus.scala 88:71]
      reqLastBeat_count_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (_reqReg_T) begin // @[Bus.scala 90:34]
      reqLastBeat_count_value <= _reqLastBeat_value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      respLastBeat_count_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (respLastBeat_fireLastBeat | _respLastBeat_fireLastBeat_T & io_resp_bits_opcode == 3'h0) begin // @[Bus.scala 99:79]
      respLastBeat_count_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (_respLastBeat_fireLastBeat_T) begin // @[Bus.scala 101:35]
      respLastBeat_count_value <= _respLastBeat_value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      beatCount_count_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (beatCount_fireLastBeat | _respLastBeat_fireLastBeat_T & io_resp_bits_opcode == 3'h0) begin // @[Bus.scala 99:79]
      beatCount_count_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (_respLastBeat_fireLastBeat_T) begin // @[Bus.scala 101:35]
      beatCount_count_value <= _beatCount_value_T_1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 131072; initvar = initvar+1)
    mem[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_rdata_addr_pipe_0 = _RAND_2[16:0];
  _RAND_3 = {1{`RANDOM}};
  reqReg_opcode = _RAND_3[2:0];
  _RAND_4 = {4{`RANDOM}};
  reqReg_size = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  reqReg_address = _RAND_5[31:0];
  _RAND_6 = {4{`RANDOM}};
  reqReg_data = _RAND_6[127:0];
  _RAND_7 = {1{`RANDOM}};
  busy = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reqLastBeat_count_value = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  respLastBeat_count_value = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  beatCount_count_value = _RAND_10[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  input         io_in_start,
  output [31:0] io_out_state_intRegState_regState_0,
  output [31:0] io_out_state_intRegState_regState_1,
  output [31:0] io_out_state_intRegState_regState_2,
  output [31:0] io_out_state_intRegState_regState_3,
  output [31:0] io_out_state_intRegState_regState_4,
  output [31:0] io_out_state_intRegState_regState_5,
  output [31:0] io_out_state_intRegState_regState_6,
  output [31:0] io_out_state_intRegState_regState_7,
  output [31:0] io_out_state_intRegState_regState_8,
  output [31:0] io_out_state_intRegState_regState_9,
  output [31:0] io_out_state_intRegState_regState_10,
  output [31:0] io_out_state_intRegState_regState_11,
  output [31:0] io_out_state_intRegState_regState_12,
  output [31:0] io_out_state_intRegState_regState_13,
  output [31:0] io_out_state_intRegState_regState_14,
  output [31:0] io_out_state_intRegState_regState_15,
  output [31:0] io_out_state_intRegState_regState_16,
  output [31:0] io_out_state_intRegState_regState_17,
  output [31:0] io_out_state_intRegState_regState_18,
  output [31:0] io_out_state_intRegState_regState_19,
  output [31:0] io_out_state_intRegState_regState_20,
  output [31:0] io_out_state_intRegState_regState_21,
  output [31:0] io_out_state_intRegState_regState_22,
  output [31:0] io_out_state_intRegState_regState_23,
  output [31:0] io_out_state_intRegState_regState_24,
  output [31:0] io_out_state_intRegState_regState_25,
  output [31:0] io_out_state_intRegState_regState_26,
  output [31:0] io_out_state_intRegState_regState_27,
  output [31:0] io_out_state_intRegState_regState_28,
  output [31:0] io_out_state_intRegState_regState_29,
  output [31:0] io_out_state_intRegState_regState_30,
  output [31:0] io_out_state_intRegState_regState_31,
  output        io_out_state_instState_commit,
  output [31:0] io_out_state_instState_pc,
  output [31:0] io_out_state_instState_inst,
  output [31:0] io_out_state_csrState_mcycle,
  output [31:0] io_out_state_csrState_mcycleh
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ife_clock; // @[Core.scala 56:21]
  wire  ife_reset; // @[Core.scala 56:21]
  wire  ife_io_in_start; // @[Core.scala 56:21]
  wire  ife_io_in_execute_bits_brTaken; // @[Core.scala 56:21]
  wire [31:0] ife_io_in_execute_bits_targetAddr; // @[Core.scala 56:21]
  wire  ife_io_out_ready; // @[Core.scala 56:21]
  wire  ife_io_out_valid; // @[Core.scala 56:21]
  wire [31:0] ife_io_out_bits_pcNext4; // @[Core.scala 56:21]
  wire  ife_io_out_bits_instState_commit; // @[Core.scala 56:21]
  wire [31:0] ife_io_out_bits_instState_pc; // @[Core.scala 56:21]
  wire [31:0] ife_io_out_bits_instState_inst; // @[Core.scala 56:21]
  wire  ife_io_tlbus_req_ready; // @[Core.scala 56:21]
  wire  ife_io_tlbus_req_valid; // @[Core.scala 56:21]
  wire [31:0] ife_io_tlbus_req_bits_address; // @[Core.scala 56:21]
  wire  ife_io_tlbus_resp_valid; // @[Core.scala 56:21]
  wire [2:0] ife_io_tlbus_resp_bits_opcode; // @[Core.scala 56:21]
  wire [127:0] ife_io_tlbus_resp_bits_data; // @[Core.scala 56:21]
  wire [31:0] ife_io_trapVec; // @[Core.scala 56:21]
  wire [31:0] ife_io_mepc; // @[Core.scala 56:21]
  wire  ife_io_excp_valid; // @[Core.scala 56:21]
  wire  ife_io_excp_bits_isMret; // @[Core.scala 56:21]
  wire  dec_clock; // @[Core.scala 64:21]
  wire  dec_reset; // @[Core.scala 64:21]
  wire  dec_io_in_ready; // @[Core.scala 64:21]
  wire  dec_io_in_valid; // @[Core.scala 64:21]
  wire [31:0] dec_io_in_bits_pcNext4; // @[Core.scala 64:21]
  wire  dec_io_in_bits_instState_commit; // @[Core.scala 64:21]
  wire [31:0] dec_io_in_bits_instState_pc; // @[Core.scala 64:21]
  wire [31:0] dec_io_in_bits_instState_inst; // @[Core.scala 64:21]
  wire  dec_io_out_ready; // @[Core.scala 64:21]
  wire  dec_io_out_valid; // @[Core.scala 64:21]
  wire  dec_io_out_bits_isBranch; // @[Core.scala 64:21]
  wire  dec_io_out_bits_isJump; // @[Core.scala 64:21]
  wire [1:0] dec_io_out_bits_resultSrc; // @[Core.scala 64:21]
  wire [4:0] dec_io_out_bits_lsuOp; // @[Core.scala 64:21]
  wire [3:0] dec_io_out_bits_aluOpSel; // @[Core.scala 64:21]
  wire  dec_io_out_bits_immSign; // @[Core.scala 64:21]
  wire  dec_io_out_bits_regWrEn; // @[Core.scala 64:21]
  wire  dec_io_out_bits_pcAddReg; // @[Core.scala 64:21]
  wire [31:0] dec_io_out_bits_pcNext4; // @[Core.scala 64:21]
  wire [31:0] dec_io_out_bits_aluIn1; // @[Core.scala 64:21]
  wire [31:0] dec_io_out_bits_aluIn2; // @[Core.scala 64:21]
  wire  dec_io_out_bits_aluIn1IsReg; // @[Core.scala 64:21]
  wire  dec_io_out_bits_aluIn2IsReg; // @[Core.scala 64:21]
  wire [31:0] dec_io_out_bits_imm; // @[Core.scala 64:21]
  wire [31:0] dec_io_out_bits_data2; // @[Core.scala 64:21]
  wire [3:0] dec_io_out_bits_excType; // @[Core.scala 64:21]
  wire [2:0] dec_io_out_bits_csrOp; // @[Core.scala 64:21]
  wire  dec_io_out_bits_instState_commit; // @[Core.scala 64:21]
  wire [31:0] dec_io_out_bits_instState_pc; // @[Core.scala 64:21]
  wire [31:0] dec_io_out_bits_instState_inst; // @[Core.scala 64:21]
  wire [4:0] dec_io_hazard_out_rs1; // @[Core.scala 64:21]
  wire [4:0] dec_io_hazard_out_rs2; // @[Core.scala 64:21]
  wire  dec_io_hazard_in_stall; // @[Core.scala 64:21]
  wire [4:0] dec_io_regfile_rs1; // @[Core.scala 64:21]
  wire [4:0] dec_io_regfile_rs2; // @[Core.scala 64:21]
  wire [31:0] dec_io_regfile_rdata1; // @[Core.scala 64:21]
  wire [31:0] dec_io_regfile_rdata2; // @[Core.scala 64:21]
  wire  dec_io_ctrl_flush; // @[Core.scala 64:21]
  wire  exe_clock; // @[Core.scala 69:21]
  wire  exe_reset; // @[Core.scala 69:21]
  wire  exe_io_in_ready; // @[Core.scala 69:21]
  wire  exe_io_in_valid; // @[Core.scala 69:21]
  wire  exe_io_in_bits_isBranch; // @[Core.scala 69:21]
  wire  exe_io_in_bits_isJump; // @[Core.scala 69:21]
  wire [1:0] exe_io_in_bits_resultSrc; // @[Core.scala 69:21]
  wire [4:0] exe_io_in_bits_lsuOp; // @[Core.scala 69:21]
  wire [3:0] exe_io_in_bits_aluOpSel; // @[Core.scala 69:21]
  wire  exe_io_in_bits_immSign; // @[Core.scala 69:21]
  wire  exe_io_in_bits_regWrEn; // @[Core.scala 69:21]
  wire  exe_io_in_bits_pcAddReg; // @[Core.scala 69:21]
  wire [31:0] exe_io_in_bits_pcNext4; // @[Core.scala 69:21]
  wire [31:0] exe_io_in_bits_aluIn1; // @[Core.scala 69:21]
  wire [31:0] exe_io_in_bits_aluIn2; // @[Core.scala 69:21]
  wire  exe_io_in_bits_aluIn1IsReg; // @[Core.scala 69:21]
  wire  exe_io_in_bits_aluIn2IsReg; // @[Core.scala 69:21]
  wire [31:0] exe_io_in_bits_imm; // @[Core.scala 69:21]
  wire [31:0] exe_io_in_bits_data2; // @[Core.scala 69:21]
  wire [3:0] exe_io_in_bits_excType; // @[Core.scala 69:21]
  wire [2:0] exe_io_in_bits_csrOp; // @[Core.scala 69:21]
  wire  exe_io_in_bits_instState_commit; // @[Core.scala 69:21]
  wire [31:0] exe_io_in_bits_instState_pc; // @[Core.scala 69:21]
  wire [31:0] exe_io_in_bits_instState_inst; // @[Core.scala 69:21]
  wire  exe_io_out_memory_ready; // @[Core.scala 69:21]
  wire  exe_io_out_memory_valid; // @[Core.scala 69:21]
  wire [1:0] exe_io_out_memory_bits_resultSrc; // @[Core.scala 69:21]
  wire [4:0] exe_io_out_memory_bits_lsuOp; // @[Core.scala 69:21]
  wire  exe_io_out_memory_bits_regWrEn; // @[Core.scala 69:21]
  wire [31:0] exe_io_out_memory_bits_aluOut; // @[Core.scala 69:21]
  wire [31:0] exe_io_out_memory_bits_data2; // @[Core.scala 69:21]
  wire [31:0] exe_io_out_memory_bits_pcNext4; // @[Core.scala 69:21]
  wire [2:0] exe_io_out_memory_bits_csrOp; // @[Core.scala 69:21]
  wire  exe_io_out_memory_bits_csrWrEn; // @[Core.scala 69:21]
  wire  exe_io_out_memory_bits_csrValid; // @[Core.scala 69:21]
  wire [31:0] exe_io_out_memory_bits_csrRdData; // @[Core.scala 69:21]
  wire [31:0] exe_io_out_memory_bits_csrWrData; // @[Core.scala 69:21]
  wire [31:0] exe_io_out_memory_bits_csrAddr; // @[Core.scala 69:21]
  wire [3:0] exe_io_out_memory_bits_excType; // @[Core.scala 69:21]
  wire  exe_io_out_memory_bits_instState_commit; // @[Core.scala 69:21]
  wire [31:0] exe_io_out_memory_bits_instState_pc; // @[Core.scala 69:21]
  wire [31:0] exe_io_out_memory_bits_instState_inst; // @[Core.scala 69:21]
  wire  exe_io_out_fetch_bits_brTaken; // @[Core.scala 69:21]
  wire [31:0] exe_io_out_fetch_bits_targetAddr; // @[Core.scala 69:21]
  wire [4:0] exe_io_hazard_out_rs1; // @[Core.scala 69:21]
  wire [4:0] exe_io_hazard_out_rs2; // @[Core.scala 69:21]
  wire [1:0] exe_io_hazard_out_resultSrc; // @[Core.scala 69:21]
  wire [4:0] exe_io_hazard_out_rd; // @[Core.scala 69:21]
  wire [1:0] exe_io_hazard_in_aluSrc1; // @[Core.scala 69:21]
  wire [1:0] exe_io_hazard_in_aluSrc2; // @[Core.scala 69:21]
  wire [31:0] exe_io_hazard_in_rdValM; // @[Core.scala 69:21]
  wire [31:0] exe_io_hazard_in_rdValW; // @[Core.scala 69:21]
  wire  exe_io_ctrl_flush; // @[Core.scala 69:21]
  wire [2:0] exe_io_csrRead_op; // @[Core.scala 69:21]
  wire  exe_io_csrRead_valid; // @[Core.scala 69:21]
  wire [11:0] exe_io_csrRead_addr; // @[Core.scala 69:21]
  wire [31:0] exe_io_csrRead_data; // @[Core.scala 69:21]
  wire  mem_clock; // @[Core.scala 74:21]
  wire  mem_reset; // @[Core.scala 74:21]
  wire  mem_io_in_ready; // @[Core.scala 74:21]
  wire [1:0] mem_io_in_bits_resultSrc; // @[Core.scala 74:21]
  wire [4:0] mem_io_in_bits_lsuOp; // @[Core.scala 74:21]
  wire  mem_io_in_bits_regWrEn; // @[Core.scala 74:21]
  wire [31:0] mem_io_in_bits_aluOut; // @[Core.scala 74:21]
  wire [31:0] mem_io_in_bits_data2; // @[Core.scala 74:21]
  wire [31:0] mem_io_in_bits_pcNext4; // @[Core.scala 74:21]
  wire [2:0] mem_io_in_bits_csrOp; // @[Core.scala 74:21]
  wire  mem_io_in_bits_csrWrEn; // @[Core.scala 74:21]
  wire  mem_io_in_bits_csrValid; // @[Core.scala 74:21]
  wire [31:0] mem_io_in_bits_csrRdData; // @[Core.scala 74:21]
  wire [31:0] mem_io_in_bits_csrWrData; // @[Core.scala 74:21]
  wire [31:0] mem_io_in_bits_csrAddr; // @[Core.scala 74:21]
  wire [3:0] mem_io_in_bits_excType; // @[Core.scala 74:21]
  wire  mem_io_in_bits_instState_commit; // @[Core.scala 74:21]
  wire [31:0] mem_io_in_bits_instState_pc; // @[Core.scala 74:21]
  wire [31:0] mem_io_in_bits_instState_inst; // @[Core.scala 74:21]
  wire  mem_io_out_ready; // @[Core.scala 74:21]
  wire  mem_io_out_valid; // @[Core.scala 74:21]
  wire [1:0] mem_io_out_bits_resultSrc; // @[Core.scala 74:21]
  wire  mem_io_out_bits_regWrEn; // @[Core.scala 74:21]
  wire [31:0] mem_io_out_bits_aluOut; // @[Core.scala 74:21]
  wire [31:0] mem_io_out_bits_pcNext4; // @[Core.scala 74:21]
  wire [2:0] mem_io_out_bits_csrOp; // @[Core.scala 74:21]
  wire  mem_io_out_bits_csrWrEn; // @[Core.scala 74:21]
  wire [31:0] mem_io_out_bits_csrRdData; // @[Core.scala 74:21]
  wire [31:0] mem_io_out_bits_csrWrData; // @[Core.scala 74:21]
  wire [11:0] mem_io_out_bits_csrAddr; // @[Core.scala 74:21]
  wire  mem_io_out_bits_instState_commit; // @[Core.scala 74:21]
  wire [31:0] mem_io_out_bits_instState_pc; // @[Core.scala 74:21]
  wire [31:0] mem_io_out_bits_instState_inst; // @[Core.scala 74:21]
  wire [31:0] mem_io_lsuData; // @[Core.scala 74:21]
  wire  mem_io_lsuOK; // @[Core.scala 74:21]
  wire  mem_io_tlbus_req_ready; // @[Core.scala 74:21]
  wire  mem_io_tlbus_req_valid; // @[Core.scala 74:21]
  wire [2:0] mem_io_tlbus_req_bits_opcode; // @[Core.scala 74:21]
  wire [31:0] mem_io_tlbus_req_bits_address; // @[Core.scala 74:21]
  wire [127:0] mem_io_tlbus_req_bits_data; // @[Core.scala 74:21]
  wire  mem_io_tlbus_resp_valid; // @[Core.scala 74:21]
  wire [2:0] mem_io_tlbus_resp_bits_opcode; // @[Core.scala 74:21]
  wire [127:0] mem_io_tlbus_resp_bits_data; // @[Core.scala 74:21]
  wire [4:0] mem_io_hazard_rd; // @[Core.scala 74:21]
  wire [31:0] mem_io_hazard_rdVal; // @[Core.scala 74:21]
  wire  mem_io_hazard_regWrEn; // @[Core.scala 74:21]
  wire  mem_io_ctrl_flush; // @[Core.scala 74:21]
  wire  mem_io_excp_valid; // @[Core.scala 74:21]
  wire  mem_io_excp_bits_isMret; // @[Core.scala 74:21]
  wire  mem_io_excp_bits_isSret; // @[Core.scala 74:21]
  wire [30:0] mem_io_excp_bits_excCause; // @[Core.scala 74:21]
  wire [31:0] mem_io_excp_bits_excPc; // @[Core.scala 74:21]
  wire  mem_io_csrBusy; // @[Core.scala 74:21]
  wire [1:0] mem_io_csrMode; // @[Core.scala 74:21]
  wire  wb_clock; // @[Core.scala 80:20]
  wire  wb_reset; // @[Core.scala 80:20]
  wire  wb_io_in_ready; // @[Core.scala 80:20]
  wire  wb_io_in_valid; // @[Core.scala 80:20]
  wire [1:0] wb_io_in_bits_resultSrc; // @[Core.scala 80:20]
  wire  wb_io_in_bits_regWrEn; // @[Core.scala 80:20]
  wire [31:0] wb_io_in_bits_aluOut; // @[Core.scala 80:20]
  wire [31:0] wb_io_in_bits_pcNext4; // @[Core.scala 80:20]
  wire [2:0] wb_io_in_bits_csrOp; // @[Core.scala 80:20]
  wire  wb_io_in_bits_csrWrEn; // @[Core.scala 80:20]
  wire [31:0] wb_io_in_bits_csrRdData; // @[Core.scala 80:20]
  wire [31:0] wb_io_in_bits_csrWrData; // @[Core.scala 80:20]
  wire [11:0] wb_io_in_bits_csrAddr; // @[Core.scala 80:20]
  wire  wb_io_in_bits_instState_commit; // @[Core.scala 80:20]
  wire [31:0] wb_io_in_bits_instState_pc; // @[Core.scala 80:20]
  wire [31:0] wb_io_in_bits_instState_inst; // @[Core.scala 80:20]
  wire  wb_io_instState_commit; // @[Core.scala 80:20]
  wire [31:0] wb_io_instState_pc; // @[Core.scala 80:20]
  wire [31:0] wb_io_instState_inst; // @[Core.scala 80:20]
  wire [4:0] wb_io_hazard_rd; // @[Core.scala 80:20]
  wire [31:0] wb_io_hazard_rdVal; // @[Core.scala 80:20]
  wire  wb_io_hazard_regWrEn; // @[Core.scala 80:20]
  wire [4:0] wb_io_regfile_rd; // @[Core.scala 80:20]
  wire  wb_io_regfile_regWrEn; // @[Core.scala 80:20]
  wire [31:0] wb_io_regfile_regWrData; // @[Core.scala 80:20]
  wire [2:0] wb_io_csrWrite_op; // @[Core.scala 80:20]
  wire [11:0] wb_io_csrWrite_addr; // @[Core.scala 80:20]
  wire [31:0] wb_io_csrWrite_data; // @[Core.scala 80:20]
  wire  wb_io_csrWrite_retired; // @[Core.scala 80:20]
  wire [31:0] wb_io_lsuData; // @[Core.scala 80:20]
  wire  pipelineCtrl_io_in_brTaken; // @[Core.scala 87:30]
  wire  pipelineCtrl_io_in_excpValid; // @[Core.scala 87:30]
  wire  pipelineCtrl_io_out_decode_flush; // @[Core.scala 87:30]
  wire  pipelineCtrl_io_out_execute_flush; // @[Core.scala 87:30]
  wire  pipelineCtrl_io_out_memory_flush; // @[Core.scala 87:30]
  wire [4:0] hazardU_io_in_decode_rs1; // @[Core.scala 97:25]
  wire [4:0] hazardU_io_in_decode_rs2; // @[Core.scala 97:25]
  wire [4:0] hazardU_io_in_execute_rs1; // @[Core.scala 97:25]
  wire [4:0] hazardU_io_in_execute_rs2; // @[Core.scala 97:25]
  wire [1:0] hazardU_io_in_execute_resultSrc; // @[Core.scala 97:25]
  wire [4:0] hazardU_io_in_execute_rd; // @[Core.scala 97:25]
  wire [4:0] hazardU_io_in_memory_rd; // @[Core.scala 97:25]
  wire [31:0] hazardU_io_in_memory_rdVal; // @[Core.scala 97:25]
  wire  hazardU_io_in_memory_regWrEn; // @[Core.scala 97:25]
  wire [4:0] hazardU_io_in_writeback_rd; // @[Core.scala 97:25]
  wire [31:0] hazardU_io_in_writeback_rdVal; // @[Core.scala 97:25]
  wire  hazardU_io_in_writeback_regWrEn; // @[Core.scala 97:25]
  wire [1:0] hazardU_io_out_execute_aluSrc1; // @[Core.scala 97:25]
  wire [1:0] hazardU_io_out_execute_aluSrc2; // @[Core.scala 97:25]
  wire [31:0] hazardU_io_out_execute_rdValM; // @[Core.scala 97:25]
  wire [31:0] hazardU_io_out_execute_rdValW; // @[Core.scala 97:25]
  wire  hazardU_io_out_decode_stall; // @[Core.scala 97:25]
  wire  regFile_clock; // @[Core.scala 106:25]
  wire  regFile_reset; // @[Core.scala 106:25]
  wire [4:0] regFile_io_r_0_addr; // @[Core.scala 106:25]
  wire [31:0] regFile_io_r_0_data; // @[Core.scala 106:25]
  wire [4:0] regFile_io_r_1_addr; // @[Core.scala 106:25]
  wire [31:0] regFile_io_r_1_data; // @[Core.scala 106:25]
  wire [4:0] regFile_io_w_0_addr; // @[Core.scala 106:25]
  wire  regFile_io_w_0_en; // @[Core.scala 106:25]
  wire [31:0] regFile_io_w_0_data; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_0; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_1; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_2; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_3; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_4; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_5; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_6; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_7; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_8; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_9; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_10; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_11; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_12; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_13; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_14; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_15; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_16; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_17; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_18; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_19; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_20; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_21; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_22; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_23; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_24; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_25; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_26; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_27; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_28; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_29; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_30; // @[Core.scala 106:25]
  wire [31:0] regFile_regState_0_regState_31; // @[Core.scala 106:25]
  wire  csrFile_clock; // @[Core.scala 118:25]
  wire  csrFile_reset; // @[Core.scala 118:25]
  wire [2:0] csrFile_io_read_op; // @[Core.scala 118:25]
  wire  csrFile_io_read_valid; // @[Core.scala 118:25]
  wire [11:0] csrFile_io_read_addr; // @[Core.scala 118:25]
  wire [31:0] csrFile_io_read_data; // @[Core.scala 118:25]
  wire [2:0] csrFile_io_write_op; // @[Core.scala 118:25]
  wire [11:0] csrFile_io_write_addr; // @[Core.scala 118:25]
  wire [31:0] csrFile_io_write_data; // @[Core.scala 118:25]
  wire  csrFile_io_write_retired; // @[Core.scala 118:25]
  wire  csrFile_io_except_valid; // @[Core.scala 118:25]
  wire  csrFile_io_except_bits_isMret; // @[Core.scala 118:25]
  wire  csrFile_io_except_bits_isSret; // @[Core.scala 118:25]
  wire [30:0] csrFile_io_except_bits_excCause; // @[Core.scala 118:25]
  wire [31:0] csrFile_io_except_bits_excPc; // @[Core.scala 118:25]
  wire [31:0] csrFile_io_except_bits_excValue; // @[Core.scala 118:25]
  wire [1:0] csrFile_io_mode; // @[Core.scala 118:25]
  wire  csrFile_io_busy; // @[Core.scala 118:25]
  wire [31:0] csrFile_io_mepc; // @[Core.scala 118:25]
  wire [31:0] csrFile_io_trapVec; // @[Core.scala 118:25]
  wire [31:0] csrFile_csrState_0_mcycle; // @[Core.scala 118:25]
  wire [31:0] csrFile_csrState_0_mcycleh; // @[Core.scala 118:25]
  wire  xbar_clock; // @[Core.scala 326:22]
  wire  xbar_reset; // @[Core.scala 326:22]
  wire  xbar_io_masterFace_in_0_ready; // @[Core.scala 326:22]
  wire  xbar_io_masterFace_in_0_valid; // @[Core.scala 326:22]
  wire [31:0] xbar_io_masterFace_in_0_bits_address; // @[Core.scala 326:22]
  wire  xbar_io_masterFace_in_1_ready; // @[Core.scala 326:22]
  wire  xbar_io_masterFace_in_1_valid; // @[Core.scala 326:22]
  wire [2:0] xbar_io_masterFace_in_1_bits_opcode; // @[Core.scala 326:22]
  wire [31:0] xbar_io_masterFace_in_1_bits_address; // @[Core.scala 326:22]
  wire [127:0] xbar_io_masterFace_in_1_bits_data; // @[Core.scala 326:22]
  wire  xbar_io_masterFace_out_0_valid; // @[Core.scala 326:22]
  wire [2:0] xbar_io_masterFace_out_0_bits_opcode; // @[Core.scala 326:22]
  wire [127:0] xbar_io_masterFace_out_0_bits_data; // @[Core.scala 326:22]
  wire  xbar_io_masterFace_out_1_valid; // @[Core.scala 326:22]
  wire [2:0] xbar_io_masterFace_out_1_bits_opcode; // @[Core.scala 326:22]
  wire [127:0] xbar_io_masterFace_out_1_bits_data; // @[Core.scala 326:22]
  wire  xbar_io_slaveFace_in_0_ready; // @[Core.scala 326:22]
  wire  xbar_io_slaveFace_in_0_valid; // @[Core.scala 326:22]
  wire [2:0] xbar_io_slaveFace_in_0_bits_opcode; // @[Core.scala 326:22]
  wire [127:0] xbar_io_slaveFace_in_0_bits_size; // @[Core.scala 326:22]
  wire [31:0] xbar_io_slaveFace_in_0_bits_address; // @[Core.scala 326:22]
  wire [127:0] xbar_io_slaveFace_in_0_bits_data; // @[Core.scala 326:22]
  wire  xbar_io_slaveFace_out_0_ready; // @[Core.scala 326:22]
  wire  xbar_io_slaveFace_out_0_valid; // @[Core.scala 326:22]
  wire [2:0] xbar_io_slaveFace_out_0_bits_opcode; // @[Core.scala 326:22]
  wire [127:0] xbar_io_slaveFace_out_0_bits_data; // @[Core.scala 326:22]
  wire  rom_clock; // @[Core.scala 327:21]
  wire  rom_reset; // @[Core.scala 327:21]
  wire  rom_io_req_ready; // @[Core.scala 327:21]
  wire  rom_io_req_valid; // @[Core.scala 327:21]
  wire [2:0] rom_io_req_bits_opcode; // @[Core.scala 327:21]
  wire [127:0] rom_io_req_bits_size; // @[Core.scala 327:21]
  wire [31:0] rom_io_req_bits_address; // @[Core.scala 327:21]
  wire [127:0] rom_io_req_bits_data; // @[Core.scala 327:21]
  wire  rom_io_resp_ready; // @[Core.scala 327:21]
  wire  rom_io_resp_valid; // @[Core.scala 327:21]
  wire [2:0] rom_io_resp_bits_opcode; // @[Core.scala 327:21]
  wire [127:0] rom_io_resp_bits_size; // @[Core.scala 327:21]
  wire [127:0] rom_io_resp_bits_data; // @[Core.scala 327:21]
  wire  ram_clock; // @[Core.scala 328:21]
  wire  ram_reset; // @[Core.scala 328:21]
  wire  ram_io_req_ready; // @[Core.scala 328:21]
  wire  ram_io_req_valid; // @[Core.scala 328:21]
  wire [2:0] ram_io_req_bits_opcode; // @[Core.scala 328:21]
  wire [127:0] ram_io_req_bits_size; // @[Core.scala 328:21]
  wire [31:0] ram_io_req_bits_address; // @[Core.scala 328:21]
  wire [127:0] ram_io_req_bits_data; // @[Core.scala 328:21]
  wire  ram_io_resp_ready; // @[Core.scala 328:21]
  wire  ram_io_resp_valid; // @[Core.scala 328:21]
  wire [2:0] ram_io_resp_bits_opcode; // @[Core.scala 328:21]
  wire [127:0] ram_io_resp_bits_size; // @[Core.scala 328:21]
  wire [127:0] ram_io_resp_bits_data; // @[Core.scala 328:21]
  reg  ife_io_in_start_REG; // @[Core.scala 57:31]
  reg  io_out_state_instState_REG_commit; // @[Core.scala 136:38]
  reg [31:0] io_out_state_instState_REG_pc; // @[Core.scala 136:38]
  reg [31:0] io_out_state_instState_REG_inst; // @[Core.scala 136:38]
  Fetch_1 ife ( // @[Core.scala 56:21]
    .clock(ife_clock),
    .reset(ife_reset),
    .io_in_start(ife_io_in_start),
    .io_in_execute_bits_brTaken(ife_io_in_execute_bits_brTaken),
    .io_in_execute_bits_targetAddr(ife_io_in_execute_bits_targetAddr),
    .io_out_ready(ife_io_out_ready),
    .io_out_valid(ife_io_out_valid),
    .io_out_bits_pcNext4(ife_io_out_bits_pcNext4),
    .io_out_bits_instState_commit(ife_io_out_bits_instState_commit),
    .io_out_bits_instState_pc(ife_io_out_bits_instState_pc),
    .io_out_bits_instState_inst(ife_io_out_bits_instState_inst),
    .io_tlbus_req_ready(ife_io_tlbus_req_ready),
    .io_tlbus_req_valid(ife_io_tlbus_req_valid),
    .io_tlbus_req_bits_address(ife_io_tlbus_req_bits_address),
    .io_tlbus_resp_valid(ife_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(ife_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(ife_io_tlbus_resp_bits_data),
    .io_trapVec(ife_io_trapVec),
    .io_mepc(ife_io_mepc),
    .io_excp_valid(ife_io_excp_valid),
    .io_excp_bits_isMret(ife_io_excp_bits_isMret)
  );
  Decode dec ( // @[Core.scala 64:21]
    .clock(dec_clock),
    .reset(dec_reset),
    .io_in_ready(dec_io_in_ready),
    .io_in_valid(dec_io_in_valid),
    .io_in_bits_pcNext4(dec_io_in_bits_pcNext4),
    .io_in_bits_instState_commit(dec_io_in_bits_instState_commit),
    .io_in_bits_instState_pc(dec_io_in_bits_instState_pc),
    .io_in_bits_instState_inst(dec_io_in_bits_instState_inst),
    .io_out_ready(dec_io_out_ready),
    .io_out_valid(dec_io_out_valid),
    .io_out_bits_isBranch(dec_io_out_bits_isBranch),
    .io_out_bits_isJump(dec_io_out_bits_isJump),
    .io_out_bits_resultSrc(dec_io_out_bits_resultSrc),
    .io_out_bits_lsuOp(dec_io_out_bits_lsuOp),
    .io_out_bits_aluOpSel(dec_io_out_bits_aluOpSel),
    .io_out_bits_immSign(dec_io_out_bits_immSign),
    .io_out_bits_regWrEn(dec_io_out_bits_regWrEn),
    .io_out_bits_pcAddReg(dec_io_out_bits_pcAddReg),
    .io_out_bits_pcNext4(dec_io_out_bits_pcNext4),
    .io_out_bits_aluIn1(dec_io_out_bits_aluIn1),
    .io_out_bits_aluIn2(dec_io_out_bits_aluIn2),
    .io_out_bits_aluIn1IsReg(dec_io_out_bits_aluIn1IsReg),
    .io_out_bits_aluIn2IsReg(dec_io_out_bits_aluIn2IsReg),
    .io_out_bits_imm(dec_io_out_bits_imm),
    .io_out_bits_data2(dec_io_out_bits_data2),
    .io_out_bits_excType(dec_io_out_bits_excType),
    .io_out_bits_csrOp(dec_io_out_bits_csrOp),
    .io_out_bits_instState_commit(dec_io_out_bits_instState_commit),
    .io_out_bits_instState_pc(dec_io_out_bits_instState_pc),
    .io_out_bits_instState_inst(dec_io_out_bits_instState_inst),
    .io_hazard_out_rs1(dec_io_hazard_out_rs1),
    .io_hazard_out_rs2(dec_io_hazard_out_rs2),
    .io_hazard_in_stall(dec_io_hazard_in_stall),
    .io_regfile_rs1(dec_io_regfile_rs1),
    .io_regfile_rs2(dec_io_regfile_rs2),
    .io_regfile_rdata1(dec_io_regfile_rdata1),
    .io_regfile_rdata2(dec_io_regfile_rdata2),
    .io_ctrl_flush(dec_io_ctrl_flush)
  );
  Execute exe ( // @[Core.scala 69:21]
    .clock(exe_clock),
    .reset(exe_reset),
    .io_in_ready(exe_io_in_ready),
    .io_in_valid(exe_io_in_valid),
    .io_in_bits_isBranch(exe_io_in_bits_isBranch),
    .io_in_bits_isJump(exe_io_in_bits_isJump),
    .io_in_bits_resultSrc(exe_io_in_bits_resultSrc),
    .io_in_bits_lsuOp(exe_io_in_bits_lsuOp),
    .io_in_bits_aluOpSel(exe_io_in_bits_aluOpSel),
    .io_in_bits_immSign(exe_io_in_bits_immSign),
    .io_in_bits_regWrEn(exe_io_in_bits_regWrEn),
    .io_in_bits_pcAddReg(exe_io_in_bits_pcAddReg),
    .io_in_bits_pcNext4(exe_io_in_bits_pcNext4),
    .io_in_bits_aluIn1(exe_io_in_bits_aluIn1),
    .io_in_bits_aluIn2(exe_io_in_bits_aluIn2),
    .io_in_bits_aluIn1IsReg(exe_io_in_bits_aluIn1IsReg),
    .io_in_bits_aluIn2IsReg(exe_io_in_bits_aluIn2IsReg),
    .io_in_bits_imm(exe_io_in_bits_imm),
    .io_in_bits_data2(exe_io_in_bits_data2),
    .io_in_bits_excType(exe_io_in_bits_excType),
    .io_in_bits_csrOp(exe_io_in_bits_csrOp),
    .io_in_bits_instState_commit(exe_io_in_bits_instState_commit),
    .io_in_bits_instState_pc(exe_io_in_bits_instState_pc),
    .io_in_bits_instState_inst(exe_io_in_bits_instState_inst),
    .io_out_memory_ready(exe_io_out_memory_ready),
    .io_out_memory_valid(exe_io_out_memory_valid),
    .io_out_memory_bits_resultSrc(exe_io_out_memory_bits_resultSrc),
    .io_out_memory_bits_lsuOp(exe_io_out_memory_bits_lsuOp),
    .io_out_memory_bits_regWrEn(exe_io_out_memory_bits_regWrEn),
    .io_out_memory_bits_aluOut(exe_io_out_memory_bits_aluOut),
    .io_out_memory_bits_data2(exe_io_out_memory_bits_data2),
    .io_out_memory_bits_pcNext4(exe_io_out_memory_bits_pcNext4),
    .io_out_memory_bits_csrOp(exe_io_out_memory_bits_csrOp),
    .io_out_memory_bits_csrWrEn(exe_io_out_memory_bits_csrWrEn),
    .io_out_memory_bits_csrValid(exe_io_out_memory_bits_csrValid),
    .io_out_memory_bits_csrRdData(exe_io_out_memory_bits_csrRdData),
    .io_out_memory_bits_csrWrData(exe_io_out_memory_bits_csrWrData),
    .io_out_memory_bits_csrAddr(exe_io_out_memory_bits_csrAddr),
    .io_out_memory_bits_excType(exe_io_out_memory_bits_excType),
    .io_out_memory_bits_instState_commit(exe_io_out_memory_bits_instState_commit),
    .io_out_memory_bits_instState_pc(exe_io_out_memory_bits_instState_pc),
    .io_out_memory_bits_instState_inst(exe_io_out_memory_bits_instState_inst),
    .io_out_fetch_bits_brTaken(exe_io_out_fetch_bits_brTaken),
    .io_out_fetch_bits_targetAddr(exe_io_out_fetch_bits_targetAddr),
    .io_hazard_out_rs1(exe_io_hazard_out_rs1),
    .io_hazard_out_rs2(exe_io_hazard_out_rs2),
    .io_hazard_out_resultSrc(exe_io_hazard_out_resultSrc),
    .io_hazard_out_rd(exe_io_hazard_out_rd),
    .io_hazard_in_aluSrc1(exe_io_hazard_in_aluSrc1),
    .io_hazard_in_aluSrc2(exe_io_hazard_in_aluSrc2),
    .io_hazard_in_rdValM(exe_io_hazard_in_rdValM),
    .io_hazard_in_rdValW(exe_io_hazard_in_rdValW),
    .io_ctrl_flush(exe_io_ctrl_flush),
    .io_csrRead_op(exe_io_csrRead_op),
    .io_csrRead_valid(exe_io_csrRead_valid),
    .io_csrRead_addr(exe_io_csrRead_addr),
    .io_csrRead_data(exe_io_csrRead_data)
  );
  Mem mem ( // @[Core.scala 74:21]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_in_ready(mem_io_in_ready),
    .io_in_bits_resultSrc(mem_io_in_bits_resultSrc),
    .io_in_bits_lsuOp(mem_io_in_bits_lsuOp),
    .io_in_bits_regWrEn(mem_io_in_bits_regWrEn),
    .io_in_bits_aluOut(mem_io_in_bits_aluOut),
    .io_in_bits_data2(mem_io_in_bits_data2),
    .io_in_bits_pcNext4(mem_io_in_bits_pcNext4),
    .io_in_bits_csrOp(mem_io_in_bits_csrOp),
    .io_in_bits_csrWrEn(mem_io_in_bits_csrWrEn),
    .io_in_bits_csrValid(mem_io_in_bits_csrValid),
    .io_in_bits_csrRdData(mem_io_in_bits_csrRdData),
    .io_in_bits_csrWrData(mem_io_in_bits_csrWrData),
    .io_in_bits_csrAddr(mem_io_in_bits_csrAddr),
    .io_in_bits_excType(mem_io_in_bits_excType),
    .io_in_bits_instState_commit(mem_io_in_bits_instState_commit),
    .io_in_bits_instState_pc(mem_io_in_bits_instState_pc),
    .io_in_bits_instState_inst(mem_io_in_bits_instState_inst),
    .io_out_ready(mem_io_out_ready),
    .io_out_valid(mem_io_out_valid),
    .io_out_bits_resultSrc(mem_io_out_bits_resultSrc),
    .io_out_bits_regWrEn(mem_io_out_bits_regWrEn),
    .io_out_bits_aluOut(mem_io_out_bits_aluOut),
    .io_out_bits_pcNext4(mem_io_out_bits_pcNext4),
    .io_out_bits_csrOp(mem_io_out_bits_csrOp),
    .io_out_bits_csrWrEn(mem_io_out_bits_csrWrEn),
    .io_out_bits_csrRdData(mem_io_out_bits_csrRdData),
    .io_out_bits_csrWrData(mem_io_out_bits_csrWrData),
    .io_out_bits_csrAddr(mem_io_out_bits_csrAddr),
    .io_out_bits_instState_commit(mem_io_out_bits_instState_commit),
    .io_out_bits_instState_pc(mem_io_out_bits_instState_pc),
    .io_out_bits_instState_inst(mem_io_out_bits_instState_inst),
    .io_lsuData(mem_io_lsuData),
    .io_lsuOK(mem_io_lsuOK),
    .io_tlbus_req_ready(mem_io_tlbus_req_ready),
    .io_tlbus_req_valid(mem_io_tlbus_req_valid),
    .io_tlbus_req_bits_opcode(mem_io_tlbus_req_bits_opcode),
    .io_tlbus_req_bits_address(mem_io_tlbus_req_bits_address),
    .io_tlbus_req_bits_data(mem_io_tlbus_req_bits_data),
    .io_tlbus_resp_valid(mem_io_tlbus_resp_valid),
    .io_tlbus_resp_bits_opcode(mem_io_tlbus_resp_bits_opcode),
    .io_tlbus_resp_bits_data(mem_io_tlbus_resp_bits_data),
    .io_hazard_rd(mem_io_hazard_rd),
    .io_hazard_rdVal(mem_io_hazard_rdVal),
    .io_hazard_regWrEn(mem_io_hazard_regWrEn),
    .io_ctrl_flush(mem_io_ctrl_flush),
    .io_excp_valid(mem_io_excp_valid),
    .io_excp_bits_isMret(mem_io_excp_bits_isMret),
    .io_excp_bits_isSret(mem_io_excp_bits_isSret),
    .io_excp_bits_excCause(mem_io_excp_bits_excCause),
    .io_excp_bits_excPc(mem_io_excp_bits_excPc),
    .io_csrBusy(mem_io_csrBusy),
    .io_csrMode(mem_io_csrMode)
  );
  WriteBack wb ( // @[Core.scala 80:20]
    .clock(wb_clock),
    .reset(wb_reset),
    .io_in_ready(wb_io_in_ready),
    .io_in_valid(wb_io_in_valid),
    .io_in_bits_resultSrc(wb_io_in_bits_resultSrc),
    .io_in_bits_regWrEn(wb_io_in_bits_regWrEn),
    .io_in_bits_aluOut(wb_io_in_bits_aluOut),
    .io_in_bits_pcNext4(wb_io_in_bits_pcNext4),
    .io_in_bits_csrOp(wb_io_in_bits_csrOp),
    .io_in_bits_csrWrEn(wb_io_in_bits_csrWrEn),
    .io_in_bits_csrRdData(wb_io_in_bits_csrRdData),
    .io_in_bits_csrWrData(wb_io_in_bits_csrWrData),
    .io_in_bits_csrAddr(wb_io_in_bits_csrAddr),
    .io_in_bits_instState_commit(wb_io_in_bits_instState_commit),
    .io_in_bits_instState_pc(wb_io_in_bits_instState_pc),
    .io_in_bits_instState_inst(wb_io_in_bits_instState_inst),
    .io_instState_commit(wb_io_instState_commit),
    .io_instState_pc(wb_io_instState_pc),
    .io_instState_inst(wb_io_instState_inst),
    .io_hazard_rd(wb_io_hazard_rd),
    .io_hazard_rdVal(wb_io_hazard_rdVal),
    .io_hazard_regWrEn(wb_io_hazard_regWrEn),
    .io_regfile_rd(wb_io_regfile_rd),
    .io_regfile_regWrEn(wb_io_regfile_regWrEn),
    .io_regfile_regWrData(wb_io_regfile_regWrData),
    .io_csrWrite_op(wb_io_csrWrite_op),
    .io_csrWrite_addr(wb_io_csrWrite_addr),
    .io_csrWrite_data(wb_io_csrWrite_data),
    .io_csrWrite_retired(wb_io_csrWrite_retired),
    .io_lsuData(wb_io_lsuData)
  );
  PipelineCtrl pipelineCtrl ( // @[Core.scala 87:30]
    .io_in_brTaken(pipelineCtrl_io_in_brTaken),
    .io_in_excpValid(pipelineCtrl_io_in_excpValid),
    .io_out_decode_flush(pipelineCtrl_io_out_decode_flush),
    .io_out_execute_flush(pipelineCtrl_io_out_execute_flush),
    .io_out_memory_flush(pipelineCtrl_io_out_memory_flush)
  );
  HazardUnit hazardU ( // @[Core.scala 97:25]
    .io_in_decode_rs1(hazardU_io_in_decode_rs1),
    .io_in_decode_rs2(hazardU_io_in_decode_rs2),
    .io_in_execute_rs1(hazardU_io_in_execute_rs1),
    .io_in_execute_rs2(hazardU_io_in_execute_rs2),
    .io_in_execute_resultSrc(hazardU_io_in_execute_resultSrc),
    .io_in_execute_rd(hazardU_io_in_execute_rd),
    .io_in_memory_rd(hazardU_io_in_memory_rd),
    .io_in_memory_rdVal(hazardU_io_in_memory_rdVal),
    .io_in_memory_regWrEn(hazardU_io_in_memory_regWrEn),
    .io_in_writeback_rd(hazardU_io_in_writeback_rd),
    .io_in_writeback_rdVal(hazardU_io_in_writeback_rdVal),
    .io_in_writeback_regWrEn(hazardU_io_in_writeback_regWrEn),
    .io_out_execute_aluSrc1(hazardU_io_out_execute_aluSrc1),
    .io_out_execute_aluSrc2(hazardU_io_out_execute_aluSrc2),
    .io_out_execute_rdValM(hazardU_io_out_execute_rdValM),
    .io_out_execute_rdValW(hazardU_io_out_execute_rdValW),
    .io_out_decode_stall(hazardU_io_out_decode_stall)
  );
  RegFile regFile ( // @[Core.scala 106:25]
    .clock(regFile_clock),
    .reset(regFile_reset),
    .io_r_0_addr(regFile_io_r_0_addr),
    .io_r_0_data(regFile_io_r_0_data),
    .io_r_1_addr(regFile_io_r_1_addr),
    .io_r_1_data(regFile_io_r_1_data),
    .io_w_0_addr(regFile_io_w_0_addr),
    .io_w_0_en(regFile_io_w_0_en),
    .io_w_0_data(regFile_io_w_0_data),
    .regState_0_regState_0(regFile_regState_0_regState_0),
    .regState_0_regState_1(regFile_regState_0_regState_1),
    .regState_0_regState_2(regFile_regState_0_regState_2),
    .regState_0_regState_3(regFile_regState_0_regState_3),
    .regState_0_regState_4(regFile_regState_0_regState_4),
    .regState_0_regState_5(regFile_regState_0_regState_5),
    .regState_0_regState_6(regFile_regState_0_regState_6),
    .regState_0_regState_7(regFile_regState_0_regState_7),
    .regState_0_regState_8(regFile_regState_0_regState_8),
    .regState_0_regState_9(regFile_regState_0_regState_9),
    .regState_0_regState_10(regFile_regState_0_regState_10),
    .regState_0_regState_11(regFile_regState_0_regState_11),
    .regState_0_regState_12(regFile_regState_0_regState_12),
    .regState_0_regState_13(regFile_regState_0_regState_13),
    .regState_0_regState_14(regFile_regState_0_regState_14),
    .regState_0_regState_15(regFile_regState_0_regState_15),
    .regState_0_regState_16(regFile_regState_0_regState_16),
    .regState_0_regState_17(regFile_regState_0_regState_17),
    .regState_0_regState_18(regFile_regState_0_regState_18),
    .regState_0_regState_19(regFile_regState_0_regState_19),
    .regState_0_regState_20(regFile_regState_0_regState_20),
    .regState_0_regState_21(regFile_regState_0_regState_21),
    .regState_0_regState_22(regFile_regState_0_regState_22),
    .regState_0_regState_23(regFile_regState_0_regState_23),
    .regState_0_regState_24(regFile_regState_0_regState_24),
    .regState_0_regState_25(regFile_regState_0_regState_25),
    .regState_0_regState_26(regFile_regState_0_regState_26),
    .regState_0_regState_27(regFile_regState_0_regState_27),
    .regState_0_regState_28(regFile_regState_0_regState_28),
    .regState_0_regState_29(regFile_regState_0_regState_29),
    .regState_0_regState_30(regFile_regState_0_regState_30),
    .regState_0_regState_31(regFile_regState_0_regState_31)
  );
  CsrFile csrFile ( // @[Core.scala 118:25]
    .clock(csrFile_clock),
    .reset(csrFile_reset),
    .io_read_op(csrFile_io_read_op),
    .io_read_valid(csrFile_io_read_valid),
    .io_read_addr(csrFile_io_read_addr),
    .io_read_data(csrFile_io_read_data),
    .io_write_op(csrFile_io_write_op),
    .io_write_addr(csrFile_io_write_addr),
    .io_write_data(csrFile_io_write_data),
    .io_write_retired(csrFile_io_write_retired),
    .io_except_valid(csrFile_io_except_valid),
    .io_except_bits_isMret(csrFile_io_except_bits_isMret),
    .io_except_bits_isSret(csrFile_io_except_bits_isSret),
    .io_except_bits_excCause(csrFile_io_except_bits_excCause),
    .io_except_bits_excPc(csrFile_io_except_bits_excPc),
    .io_except_bits_excValue(csrFile_io_except_bits_excValue),
    .io_mode(csrFile_io_mode),
    .io_busy(csrFile_io_busy),
    .io_mepc(csrFile_io_mepc),
    .io_trapVec(csrFile_io_trapVec),
    .csrState_0_mcycle(csrFile_csrState_0_mcycle),
    .csrState_0_mcycleh(csrFile_csrState_0_mcycleh)
  );
  TLXbar xbar ( // @[Core.scala 326:22]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_masterFace_in_0_ready(xbar_io_masterFace_in_0_ready),
    .io_masterFace_in_0_valid(xbar_io_masterFace_in_0_valid),
    .io_masterFace_in_0_bits_address(xbar_io_masterFace_in_0_bits_address),
    .io_masterFace_in_1_ready(xbar_io_masterFace_in_1_ready),
    .io_masterFace_in_1_valid(xbar_io_masterFace_in_1_valid),
    .io_masterFace_in_1_bits_opcode(xbar_io_masterFace_in_1_bits_opcode),
    .io_masterFace_in_1_bits_address(xbar_io_masterFace_in_1_bits_address),
    .io_masterFace_in_1_bits_data(xbar_io_masterFace_in_1_bits_data),
    .io_masterFace_out_0_valid(xbar_io_masterFace_out_0_valid),
    .io_masterFace_out_0_bits_opcode(xbar_io_masterFace_out_0_bits_opcode),
    .io_masterFace_out_0_bits_data(xbar_io_masterFace_out_0_bits_data),
    .io_masterFace_out_1_valid(xbar_io_masterFace_out_1_valid),
    .io_masterFace_out_1_bits_opcode(xbar_io_masterFace_out_1_bits_opcode),
    .io_masterFace_out_1_bits_data(xbar_io_masterFace_out_1_bits_data),
    .io_slaveFace_in_0_ready(xbar_io_slaveFace_in_0_ready),
    .io_slaveFace_in_0_valid(xbar_io_slaveFace_in_0_valid),
    .io_slaveFace_in_0_bits_opcode(xbar_io_slaveFace_in_0_bits_opcode),
    .io_slaveFace_in_0_bits_size(xbar_io_slaveFace_in_0_bits_size),
    .io_slaveFace_in_0_bits_address(xbar_io_slaveFace_in_0_bits_address),
    .io_slaveFace_in_0_bits_data(xbar_io_slaveFace_in_0_bits_data),
    .io_slaveFace_out_0_ready(xbar_io_slaveFace_out_0_ready),
    .io_slaveFace_out_0_valid(xbar_io_slaveFace_out_0_valid),
    .io_slaveFace_out_0_bits_opcode(xbar_io_slaveFace_out_0_bits_opcode),
    .io_slaveFace_out_0_bits_data(xbar_io_slaveFace_out_0_bits_data)
  );
  SingleROM rom ( // @[Core.scala 327:21]
    .clock(rom_clock),
    .reset(rom_reset),
    .io_req_ready(rom_io_req_ready),
    .io_req_valid(rom_io_req_valid),
    .io_req_bits_opcode(rom_io_req_bits_opcode),
    .io_req_bits_size(rom_io_req_bits_size),
    .io_req_bits_address(rom_io_req_bits_address),
    .io_req_bits_data(rom_io_req_bits_data),
    .io_resp_ready(rom_io_resp_ready),
    .io_resp_valid(rom_io_resp_valid),
    .io_resp_bits_opcode(rom_io_resp_bits_opcode),
    .io_resp_bits_size(rom_io_resp_bits_size),
    .io_resp_bits_data(rom_io_resp_bits_data)
  );
  SingleROM ram ( // @[Core.scala 328:21]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_req_ready(ram_io_req_ready),
    .io_req_valid(ram_io_req_valid),
    .io_req_bits_opcode(ram_io_req_bits_opcode),
    .io_req_bits_size(ram_io_req_bits_size),
    .io_req_bits_address(ram_io_req_bits_address),
    .io_req_bits_data(ram_io_req_bits_data),
    .io_resp_ready(ram_io_resp_ready),
    .io_resp_valid(ram_io_resp_valid),
    .io_resp_bits_opcode(ram_io_resp_bits_opcode),
    .io_resp_bits_size(ram_io_resp_bits_size),
    .io_resp_bits_data(ram_io_resp_bits_data)
  );
  assign io_out_state_intRegState_regState_0 = regFile_regState_0_regState_0; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_1 = regFile_regState_0_regState_1; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_2 = regFile_regState_0_regState_2; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_3 = regFile_regState_0_regState_3; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_4 = regFile_regState_0_regState_4; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_5 = regFile_regState_0_regState_5; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_6 = regFile_regState_0_regState_6; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_7 = regFile_regState_0_regState_7; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_8 = regFile_regState_0_regState_8; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_9 = regFile_regState_0_regState_9; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_10 = regFile_regState_0_regState_10; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_11 = regFile_regState_0_regState_11; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_12 = regFile_regState_0_regState_12; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_13 = regFile_regState_0_regState_13; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_14 = regFile_regState_0_regState_14; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_15 = regFile_regState_0_regState_15; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_16 = regFile_regState_0_regState_16; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_17 = regFile_regState_0_regState_17; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_18 = regFile_regState_0_regState_18; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_19 = regFile_regState_0_regState_19; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_20 = regFile_regState_0_regState_20; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_21 = regFile_regState_0_regState_21; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_22 = regFile_regState_0_regState_22; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_23 = regFile_regState_0_regState_23; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_24 = regFile_regState_0_regState_24; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_25 = regFile_regState_0_regState_25; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_26 = regFile_regState_0_regState_26; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_27 = regFile_regState_0_regState_27; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_28 = regFile_regState_0_regState_28; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_29 = regFile_regState_0_regState_29; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_30 = regFile_regState_0_regState_30; // @[Core.scala 130:28]
  assign io_out_state_intRegState_regState_31 = regFile_regState_0_regState_31; // @[Core.scala 130:28]
  assign io_out_state_instState_commit = io_out_state_instState_REG_commit; // @[Core.scala 136:28]
  assign io_out_state_instState_pc = io_out_state_instState_REG_pc; // @[Core.scala 136:28]
  assign io_out_state_instState_inst = io_out_state_instState_REG_inst; // @[Core.scala 136:28]
  assign io_out_state_csrState_mcycle = csrFile_csrState_0_mcycle; // @[Core.scala 133:28]
  assign io_out_state_csrState_mcycleh = csrFile_csrState_0_mcycleh; // @[Core.scala 133:28]
  assign ife_clock = clock;
  assign ife_reset = reset;
  assign ife_io_in_start = ife_io_in_start_REG; // @[Core.scala 57:21]
  assign ife_io_in_execute_bits_brTaken = exe_io_out_fetch_bits_brTaken; // @[Core.scala 71:23]
  assign ife_io_in_execute_bits_targetAddr = exe_io_out_fetch_bits_targetAddr; // @[Core.scala 71:23]
  assign ife_io_out_ready = dec_io_in_ready; // @[Core.scala 65:15]
  assign ife_io_tlbus_req_ready = xbar_io_masterFace_in_0_ready; // @[Core.scala 332:22]
  assign ife_io_tlbus_resp_valid = xbar_io_masterFace_out_0_valid; // @[Core.scala 333:23]
  assign ife_io_tlbus_resp_bits_opcode = xbar_io_masterFace_out_0_bits_opcode; // @[Core.scala 333:23]
  assign ife_io_tlbus_resp_bits_data = xbar_io_masterFace_out_0_bits_data; // @[Core.scala 333:23]
  assign ife_io_trapVec = csrFile_io_trapVec; // @[Core.scala 125:13 51:23]
  assign ife_io_mepc = csrFile_io_mepc; // @[Core.scala 126:10 52:20]
  assign ife_io_excp_valid = mem_io_excp_valid; // @[Core.scala 77:17]
  assign ife_io_excp_bits_isMret = mem_io_excp_bits_isMret; // @[Core.scala 77:17]
  assign dec_clock = clock;
  assign dec_reset = reset;
  assign dec_io_in_valid = ife_io_out_valid; // @[Core.scala 65:15]
  assign dec_io_in_bits_pcNext4 = ife_io_out_bits_pcNext4; // @[Core.scala 65:15]
  assign dec_io_in_bits_instState_commit = ife_io_out_bits_instState_commit; // @[Core.scala 65:15]
  assign dec_io_in_bits_instState_pc = ife_io_out_bits_instState_pc; // @[Core.scala 65:15]
  assign dec_io_in_bits_instState_inst = ife_io_out_bits_instState_inst; // @[Core.scala 65:15]
  assign dec_io_out_ready = exe_io_in_ready; // @[Core.scala 70:15]
  assign dec_io_hazard_in_stall = hazardU_io_out_decode_stall; // @[Core.scala 103:14 49:24]
  assign dec_io_regfile_rdata1 = regFile_io_r_0_data; // @[Core.scala 111:27]
  assign dec_io_regfile_rdata2 = regFile_io_r_1_data; // @[Core.scala 112:27]
  assign dec_io_ctrl_flush = pipelineCtrl_io_out_decode_flush; // @[Core.scala 91:17]
  assign exe_clock = clock;
  assign exe_reset = reset;
  assign exe_io_in_valid = dec_io_out_valid; // @[Core.scala 70:15]
  assign exe_io_in_bits_isBranch = dec_io_out_bits_isBranch; // @[Core.scala 70:15]
  assign exe_io_in_bits_isJump = dec_io_out_bits_isJump; // @[Core.scala 70:15]
  assign exe_io_in_bits_resultSrc = dec_io_out_bits_resultSrc; // @[Core.scala 70:15]
  assign exe_io_in_bits_lsuOp = dec_io_out_bits_lsuOp; // @[Core.scala 70:15]
  assign exe_io_in_bits_aluOpSel = dec_io_out_bits_aluOpSel; // @[Core.scala 70:15]
  assign exe_io_in_bits_immSign = dec_io_out_bits_immSign; // @[Core.scala 70:15]
  assign exe_io_in_bits_regWrEn = dec_io_out_bits_regWrEn; // @[Core.scala 70:15]
  assign exe_io_in_bits_pcAddReg = dec_io_out_bits_pcAddReg; // @[Core.scala 70:15]
  assign exe_io_in_bits_pcNext4 = dec_io_out_bits_pcNext4; // @[Core.scala 70:15]
  assign exe_io_in_bits_aluIn1 = dec_io_out_bits_aluIn1; // @[Core.scala 70:15]
  assign exe_io_in_bits_aluIn2 = dec_io_out_bits_aluIn2; // @[Core.scala 70:15]
  assign exe_io_in_bits_aluIn1IsReg = dec_io_out_bits_aluIn1IsReg; // @[Core.scala 70:15]
  assign exe_io_in_bits_aluIn2IsReg = dec_io_out_bits_aluIn2IsReg; // @[Core.scala 70:15]
  assign exe_io_in_bits_imm = dec_io_out_bits_imm; // @[Core.scala 70:15]
  assign exe_io_in_bits_data2 = dec_io_out_bits_data2; // @[Core.scala 70:15]
  assign exe_io_in_bits_excType = dec_io_out_bits_excType; // @[Core.scala 70:15]
  assign exe_io_in_bits_csrOp = dec_io_out_bits_csrOp; // @[Core.scala 70:15]
  assign exe_io_in_bits_instState_commit = dec_io_out_bits_instState_commit; // @[Core.scala 70:15]
  assign exe_io_in_bits_instState_pc = dec_io_out_bits_instState_pc; // @[Core.scala 70:15]
  assign exe_io_in_bits_instState_inst = dec_io_out_bits_instState_inst; // @[Core.scala 70:15]
  assign exe_io_out_memory_ready = mem_io_in_ready; // @[Core.scala 75:15]
  assign exe_io_hazard_in_aluSrc1 = hazardU_io_out_execute_aluSrc1; // @[Core.scala 102:29]
  assign exe_io_hazard_in_aluSrc2 = hazardU_io_out_execute_aluSrc2; // @[Core.scala 102:29]
  assign exe_io_hazard_in_rdValM = hazardU_io_out_execute_rdValM; // @[Core.scala 102:29]
  assign exe_io_hazard_in_rdValW = hazardU_io_out_execute_rdValW; // @[Core.scala 102:29]
  assign exe_io_ctrl_flush = pipelineCtrl_io_out_execute_flush; // @[Core.scala 92:17]
  assign exe_io_csrRead_valid = csrFile_io_read_valid; // @[Core.scala 121:21]
  assign exe_io_csrRead_data = csrFile_io_read_data; // @[Core.scala 121:21]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_in_bits_resultSrc = exe_io_out_memory_bits_resultSrc; // @[Core.scala 75:15]
  assign mem_io_in_bits_lsuOp = exe_io_out_memory_bits_lsuOp; // @[Core.scala 75:15]
  assign mem_io_in_bits_regWrEn = exe_io_out_memory_bits_regWrEn; // @[Core.scala 75:15]
  assign mem_io_in_bits_aluOut = exe_io_out_memory_bits_aluOut; // @[Core.scala 75:15]
  assign mem_io_in_bits_data2 = exe_io_out_memory_bits_data2; // @[Core.scala 75:15]
  assign mem_io_in_bits_pcNext4 = exe_io_out_memory_bits_pcNext4; // @[Core.scala 75:15]
  assign mem_io_in_bits_csrOp = exe_io_out_memory_bits_csrOp; // @[Core.scala 75:15]
  assign mem_io_in_bits_csrWrEn = exe_io_out_memory_bits_csrWrEn; // @[Core.scala 75:15]
  assign mem_io_in_bits_csrValid = exe_io_out_memory_bits_csrValid; // @[Core.scala 75:15]
  assign mem_io_in_bits_csrRdData = exe_io_out_memory_bits_csrRdData; // @[Core.scala 75:15]
  assign mem_io_in_bits_csrWrData = exe_io_out_memory_bits_csrWrData; // @[Core.scala 75:15]
  assign mem_io_in_bits_csrAddr = exe_io_out_memory_bits_csrAddr; // @[Core.scala 75:15]
  assign mem_io_in_bits_excType = exe_io_out_memory_bits_excType; // @[Core.scala 75:15]
  assign mem_io_in_bits_instState_commit = exe_io_out_memory_bits_instState_commit; // @[Core.scala 75:15]
  assign mem_io_in_bits_instState_pc = exe_io_out_memory_bits_instState_pc; // @[Core.scala 75:15]
  assign mem_io_in_bits_instState_inst = exe_io_out_memory_bits_instState_inst; // @[Core.scala 75:15]
  assign mem_io_out_ready = wb_io_in_ready; // @[Core.scala 81:14]
  assign mem_io_tlbus_req_ready = xbar_io_masterFace_in_1_ready; // @[Core.scala 335:22]
  assign mem_io_tlbus_resp_valid = xbar_io_masterFace_out_1_valid; // @[Core.scala 336:23]
  assign mem_io_tlbus_resp_bits_opcode = xbar_io_masterFace_out_1_bits_opcode; // @[Core.scala 336:23]
  assign mem_io_tlbus_resp_bits_data = xbar_io_masterFace_out_1_bits_data; // @[Core.scala 336:23]
  assign mem_io_ctrl_flush = pipelineCtrl_io_out_memory_flush; // @[Core.scala 93:17]
  assign mem_io_csrBusy = csrFile_io_busy; // @[Core.scala 123:20]
  assign mem_io_csrMode = csrFile_io_mode; // @[Core.scala 124:20]
  assign wb_clock = clock;
  assign wb_reset = reset;
  assign wb_io_in_valid = mem_io_out_valid; // @[Core.scala 81:14]
  assign wb_io_in_bits_resultSrc = mem_io_out_bits_resultSrc; // @[Core.scala 81:14]
  assign wb_io_in_bits_regWrEn = mem_io_out_bits_regWrEn; // @[Core.scala 81:14]
  assign wb_io_in_bits_aluOut = mem_io_out_bits_aluOut; // @[Core.scala 81:14]
  assign wb_io_in_bits_pcNext4 = mem_io_out_bits_pcNext4; // @[Core.scala 81:14]
  assign wb_io_in_bits_csrOp = mem_io_out_bits_csrOp; // @[Core.scala 81:14]
  assign wb_io_in_bits_csrWrEn = mem_io_out_bits_csrWrEn; // @[Core.scala 81:14]
  assign wb_io_in_bits_csrRdData = mem_io_out_bits_csrRdData; // @[Core.scala 81:14]
  assign wb_io_in_bits_csrWrData = mem_io_out_bits_csrWrData; // @[Core.scala 81:14]
  assign wb_io_in_bits_csrAddr = mem_io_out_bits_csrAddr; // @[Core.scala 81:14]
  assign wb_io_in_bits_instState_commit = mem_io_out_bits_instState_commit; // @[Core.scala 81:14]
  assign wb_io_in_bits_instState_pc = mem_io_out_bits_instState_pc; // @[Core.scala 81:14]
  assign wb_io_in_bits_instState_inst = mem_io_out_bits_instState_inst; // @[Core.scala 81:14]
  assign wb_io_lsuData = mem_io_lsuData; // @[Core.scala 82:19]
  assign pipelineCtrl_io_in_brTaken = exe_io_out_fetch_bits_brTaken; // @[Core.scala 89:34]
  assign pipelineCtrl_io_in_excpValid = mem_io_excp_valid; // @[Core.scala 88:34]
  assign hazardU_io_in_decode_rs1 = dec_io_hazard_out_rs1; // @[Core.scala 98:29]
  assign hazardU_io_in_decode_rs2 = dec_io_hazard_out_rs2; // @[Core.scala 98:29]
  assign hazardU_io_in_execute_rs1 = exe_io_hazard_out_rs1; // @[Core.scala 99:29]
  assign hazardU_io_in_execute_rs2 = exe_io_hazard_out_rs2; // @[Core.scala 99:29]
  assign hazardU_io_in_execute_resultSrc = exe_io_hazard_out_resultSrc; // @[Core.scala 99:29]
  assign hazardU_io_in_execute_rd = exe_io_hazard_out_rd; // @[Core.scala 99:29]
  assign hazardU_io_in_memory_rd = mem_io_hazard_rd; // @[Core.scala 100:29]
  assign hazardU_io_in_memory_rdVal = mem_io_hazard_rdVal; // @[Core.scala 100:29]
  assign hazardU_io_in_memory_regWrEn = mem_io_hazard_regWrEn; // @[Core.scala 100:29]
  assign hazardU_io_in_writeback_rd = wb_io_hazard_rd; // @[Core.scala 101:29]
  assign hazardU_io_in_writeback_rdVal = wb_io_hazard_rdVal; // @[Core.scala 101:29]
  assign hazardU_io_in_writeback_regWrEn = wb_io_hazard_regWrEn; // @[Core.scala 101:29]
  assign regFile_clock = clock;
  assign regFile_reset = reset;
  assign regFile_io_r_0_addr = dec_io_regfile_rs1; // @[Core.scala 109:26]
  assign regFile_io_r_1_addr = dec_io_regfile_rs2; // @[Core.scala 110:26]
  assign regFile_io_w_0_addr = wb_io_regfile_rd; // @[Core.scala 114:26]
  assign regFile_io_w_0_en = wb_io_regfile_regWrEn; // @[Core.scala 113:24]
  assign regFile_io_w_0_data = wb_io_regfile_regWrData; // @[Core.scala 115:26]
  assign csrFile_clock = clock;
  assign csrFile_reset = reset;
  assign csrFile_io_read_op = exe_io_csrRead_op; // @[Core.scala 121:21]
  assign csrFile_io_read_addr = exe_io_csrRead_addr; // @[Core.scala 121:21]
  assign csrFile_io_write_op = wb_io_csrWrite_op; // @[Core.scala 122:22]
  assign csrFile_io_write_addr = wb_io_csrWrite_addr; // @[Core.scala 122:22]
  assign csrFile_io_write_data = wb_io_csrWrite_data; // @[Core.scala 122:22]
  assign csrFile_io_write_retired = wb_io_csrWrite_retired; // @[Core.scala 122:22]
  assign csrFile_io_except_valid = mem_io_excp_valid; // @[Core.scala 120:23]
  assign csrFile_io_except_bits_isMret = mem_io_excp_bits_isMret; // @[Core.scala 120:23]
  assign csrFile_io_except_bits_isSret = mem_io_excp_bits_isSret; // @[Core.scala 120:23]
  assign csrFile_io_except_bits_excCause = mem_io_excp_bits_excCause; // @[Core.scala 120:23]
  assign csrFile_io_except_bits_excPc = mem_io_excp_bits_excPc; // @[Core.scala 120:23]
  assign csrFile_io_except_bits_excValue = 32'h0; // @[Core.scala 120:23]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_masterFace_in_0_valid = ife_io_tlbus_req_valid; // @[Core.scala 332:22]
  assign xbar_io_masterFace_in_0_bits_address = ife_io_tlbus_req_bits_address; // @[Core.scala 332:22]
  assign xbar_io_masterFace_in_1_valid = mem_io_tlbus_req_valid; // @[Core.scala 335:22]
  assign xbar_io_masterFace_in_1_bits_opcode = mem_io_tlbus_req_bits_opcode; // @[Core.scala 335:22]
  assign xbar_io_masterFace_in_1_bits_address = mem_io_tlbus_req_bits_address; // @[Core.scala 335:22]
  assign xbar_io_masterFace_in_1_bits_data = mem_io_tlbus_req_bits_data; // @[Core.scala 335:22]
  assign xbar_io_slaveFace_in_0_ready = rom_io_req_ready; // @[Core.scala 340:16]
  assign xbar_io_slaveFace_out_0_valid = rom_io_resp_valid; // @[Core.scala 341:17]
  assign xbar_io_slaveFace_out_0_bits_opcode = rom_io_resp_bits_opcode; // @[Core.scala 341:17]
  assign xbar_io_slaveFace_out_0_bits_data = rom_io_resp_bits_data; // @[Core.scala 341:17]
  assign rom_clock = clock;
  assign rom_reset = reset;
  assign rom_io_req_valid = xbar_io_slaveFace_in_0_valid; // @[Core.scala 340:16]
  assign rom_io_req_bits_opcode = xbar_io_slaveFace_in_0_bits_opcode; // @[Core.scala 340:16]
  assign rom_io_req_bits_size = xbar_io_slaveFace_in_0_bits_size; // @[Core.scala 340:16]
  assign rom_io_req_bits_address = xbar_io_slaveFace_in_0_bits_address; // @[Core.scala 340:16]
  assign rom_io_req_bits_data = xbar_io_slaveFace_in_0_bits_data; // @[Core.scala 340:16]
  assign rom_io_resp_ready = xbar_io_slaveFace_out_0_ready; // @[Core.scala 341:17]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_req_valid = 1'h0;
  assign ram_io_req_bits_opcode = 3'h0;
  assign ram_io_req_bits_size = 128'h0;
  assign ram_io_req_bits_address = 32'h0;
  assign ram_io_req_bits_data = 128'h0;
  assign ram_io_resp_ready = 1'h0;
  always @(posedge clock) begin
    ife_io_in_start_REG <= io_in_start; // @[Core.scala 57:31]
    io_out_state_instState_REG_commit <= wb_io_instState_commit; // @[Core.scala 136:38]
    io_out_state_instState_REG_pc <= wb_io_instState_pc; // @[Core.scala 136:38]
    io_out_state_instState_REG_inst <= wb_io_instState_inst; // @[Core.scala 136:38]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ife_io_in_start_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_out_state_instState_REG_commit = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_out_state_instState_REG_pc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_out_state_instState_REG_inst = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
