module BankRAM_2P_100(
  input        clock,
  input        reset,
  input  [8:0] io_r_addr,
  output [1:0] io_r_data,
  input        io_w_en,
  input  [8:0] io_w_addr,
  input  [1:0] io_w_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] mem [0:511]; // @[SRAM_1.scala 63:26]
  wire  mem_io_r_data_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_io_r_data_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_io_r_data_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_1_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_1_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_2_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_2_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_3_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_3_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_4_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_4_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_5_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_5_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_6_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_6_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_7_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_7_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_8_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_8_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_9_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_9_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_10_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_10_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_11_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_11_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_12_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_12_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_13_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_13_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_14_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_14_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_15_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_15_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_16_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_16_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_17_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_17_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_18_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_18_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_19_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_19_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_20_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_20_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_21_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_21_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_22_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_22_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_23_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_23_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_24_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_24_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_25_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_25_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_26_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_26_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_27_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_27_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_28_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_28_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_29_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_29_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_30_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_30_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_31_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_31_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_32_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_32_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_33_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_33_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_34_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_34_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_35_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_35_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_36_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_36_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_37_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_37_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_38_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_38_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_39_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_39_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_40_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_40_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_41_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_41_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_42_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_42_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_43_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_43_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_44_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_44_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_45_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_45_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_46_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_46_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_47_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_47_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_48_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_48_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_49_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_49_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_50_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_50_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_51_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_51_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_52_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_52_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_53_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_53_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_54_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_54_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_55_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_55_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_56_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_56_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_57_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_57_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_58_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_58_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_59_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_59_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_60_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_60_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_61_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_61_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_62_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_62_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_63_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_63_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_64_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_64_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_65_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_65_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_66_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_66_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_67_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_67_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_68_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_68_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_69_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_69_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_70_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_70_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_71_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_71_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_72_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_72_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_73_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_73_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_74_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_74_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_75_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_75_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_76_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_76_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_77_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_77_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_78_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_78_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_79_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_79_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_80_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_80_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_81_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_81_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_82_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_82_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_83_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_83_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_84_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_84_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_85_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_85_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_86_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_86_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_87_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_87_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_88_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_88_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_89_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_89_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_90_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_90_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_91_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_91_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_92_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_92_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_93_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_93_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_94_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_94_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_95_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_95_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_96_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_96_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_97_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_97_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_98_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_98_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_99_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_99_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_100_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_100_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_101_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_101_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_102_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_102_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_103_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_103_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_104_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_104_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_105_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_105_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_106_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_106_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_107_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_107_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_108_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_108_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_109_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_109_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_110_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_110_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_111_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_111_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_112_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_112_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_113_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_113_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_114_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_114_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_115_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_115_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_116_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_116_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_117_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_117_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_118_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_118_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_119_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_119_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_120_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_120_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_121_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_121_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_122_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_122_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_123_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_123_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_124_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_124_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_125_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_125_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_126_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_126_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_127_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_127_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_128_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_128_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_129_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_129_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_130_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_130_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_131_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_131_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_132_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_132_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_133_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_133_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_134_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_134_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_135_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_135_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_136_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_136_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_137_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_137_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_138_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_138_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_139_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_139_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_140_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_140_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_141_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_141_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_142_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_142_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_143_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_143_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_144_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_144_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_145_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_145_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_146_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_146_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_147_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_147_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_148_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_148_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_149_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_149_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_150_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_150_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_151_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_151_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_152_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_152_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_153_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_153_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_154_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_154_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_155_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_155_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_156_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_156_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_157_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_157_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_158_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_158_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_159_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_159_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_160_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_160_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_161_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_161_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_162_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_162_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_163_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_163_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_164_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_164_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_165_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_165_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_166_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_166_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_167_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_167_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_168_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_168_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_169_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_169_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_170_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_170_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_171_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_171_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_172_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_172_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_173_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_173_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_174_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_174_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_175_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_175_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_176_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_176_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_177_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_177_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_178_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_178_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_179_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_179_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_180_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_180_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_181_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_181_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_182_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_182_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_183_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_183_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_184_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_184_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_185_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_185_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_186_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_186_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_187_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_187_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_188_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_188_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_189_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_189_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_190_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_190_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_191_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_191_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_192_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_192_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_193_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_193_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_194_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_194_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_195_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_195_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_196_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_196_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_197_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_197_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_198_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_198_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_199_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_199_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_200_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_200_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_201_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_201_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_202_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_202_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_203_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_203_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_204_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_204_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_205_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_205_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_206_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_206_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_207_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_207_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_208_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_208_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_209_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_209_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_210_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_210_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_211_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_211_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_212_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_212_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_213_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_213_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_214_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_214_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_215_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_215_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_216_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_216_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_217_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_217_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_218_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_218_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_219_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_219_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_220_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_220_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_221_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_221_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_222_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_222_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_223_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_223_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_224_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_224_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_225_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_225_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_226_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_226_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_227_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_227_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_228_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_228_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_229_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_229_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_230_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_230_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_231_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_231_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_232_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_232_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_233_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_233_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_234_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_234_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_235_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_235_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_236_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_236_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_237_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_237_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_238_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_238_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_239_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_239_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_240_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_240_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_241_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_241_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_242_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_242_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_243_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_243_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_244_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_244_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_245_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_245_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_246_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_246_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_247_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_247_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_248_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_248_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_249_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_249_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_250_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_250_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_251_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_251_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_252_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_252_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_253_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_253_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_254_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_254_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_255_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_255_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_256_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_256_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_257_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_257_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_257_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_257_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_258_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_258_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_258_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_258_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_259_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_259_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_259_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_259_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_260_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_260_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_260_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_260_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_261_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_261_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_261_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_261_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_262_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_262_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_262_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_262_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_263_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_263_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_263_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_263_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_264_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_264_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_264_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_264_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_265_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_265_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_265_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_265_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_266_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_266_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_266_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_266_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_267_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_267_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_267_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_267_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_268_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_268_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_268_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_268_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_269_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_269_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_269_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_269_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_270_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_270_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_270_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_270_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_271_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_271_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_271_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_271_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_272_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_272_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_272_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_272_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_273_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_273_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_273_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_273_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_274_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_274_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_274_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_274_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_275_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_275_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_275_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_275_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_276_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_276_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_276_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_276_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_277_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_277_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_277_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_277_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_278_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_278_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_278_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_278_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_279_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_279_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_279_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_279_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_280_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_280_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_280_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_280_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_281_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_281_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_281_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_281_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_282_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_282_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_282_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_282_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_283_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_283_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_283_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_283_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_284_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_284_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_284_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_284_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_285_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_285_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_285_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_285_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_286_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_286_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_286_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_286_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_287_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_287_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_287_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_287_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_288_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_288_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_288_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_288_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_289_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_289_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_289_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_289_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_290_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_290_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_290_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_290_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_291_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_291_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_291_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_291_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_292_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_292_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_292_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_292_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_293_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_293_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_293_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_293_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_294_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_294_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_294_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_294_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_295_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_295_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_295_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_295_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_296_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_296_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_296_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_296_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_297_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_297_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_297_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_297_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_298_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_298_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_298_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_298_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_299_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_299_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_299_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_299_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_300_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_300_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_300_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_300_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_301_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_301_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_301_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_301_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_302_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_302_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_302_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_302_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_303_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_303_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_303_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_303_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_304_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_304_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_304_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_304_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_305_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_305_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_305_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_305_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_306_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_306_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_306_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_306_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_307_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_307_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_307_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_307_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_308_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_308_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_308_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_308_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_309_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_309_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_309_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_309_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_310_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_310_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_310_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_310_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_311_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_311_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_311_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_311_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_312_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_312_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_312_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_312_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_313_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_313_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_313_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_313_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_314_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_314_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_314_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_314_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_315_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_315_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_315_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_315_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_316_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_316_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_316_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_316_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_317_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_317_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_317_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_317_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_318_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_318_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_318_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_318_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_319_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_319_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_319_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_319_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_320_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_320_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_320_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_320_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_321_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_321_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_321_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_321_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_322_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_322_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_322_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_322_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_323_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_323_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_323_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_323_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_324_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_324_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_324_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_324_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_325_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_325_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_325_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_325_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_326_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_326_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_326_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_326_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_327_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_327_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_327_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_327_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_328_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_328_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_328_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_328_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_329_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_329_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_329_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_329_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_330_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_330_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_330_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_330_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_331_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_331_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_331_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_331_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_332_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_332_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_332_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_332_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_333_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_333_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_333_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_333_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_334_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_334_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_334_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_334_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_335_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_335_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_335_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_335_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_336_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_336_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_336_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_336_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_337_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_337_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_337_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_337_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_338_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_338_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_338_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_338_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_339_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_339_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_339_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_339_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_340_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_340_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_340_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_340_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_341_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_341_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_341_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_341_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_342_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_342_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_342_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_342_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_343_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_343_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_343_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_343_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_344_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_344_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_344_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_344_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_345_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_345_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_345_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_345_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_346_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_346_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_346_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_346_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_347_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_347_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_347_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_347_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_348_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_348_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_348_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_348_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_349_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_349_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_349_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_349_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_350_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_350_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_350_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_350_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_351_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_351_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_351_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_351_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_352_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_352_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_352_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_352_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_353_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_353_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_353_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_353_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_354_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_354_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_354_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_354_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_355_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_355_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_355_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_355_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_356_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_356_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_356_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_356_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_357_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_357_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_357_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_357_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_358_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_358_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_358_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_358_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_359_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_359_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_359_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_359_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_360_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_360_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_360_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_360_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_361_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_361_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_361_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_361_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_362_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_362_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_362_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_362_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_363_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_363_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_363_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_363_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_364_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_364_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_364_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_364_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_365_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_365_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_365_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_365_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_366_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_366_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_366_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_366_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_367_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_367_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_367_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_367_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_368_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_368_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_368_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_368_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_369_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_369_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_369_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_369_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_370_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_370_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_370_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_370_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_371_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_371_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_371_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_371_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_372_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_372_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_372_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_372_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_373_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_373_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_373_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_373_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_374_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_374_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_374_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_374_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_375_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_375_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_375_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_375_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_376_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_376_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_376_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_376_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_377_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_377_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_377_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_377_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_378_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_378_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_378_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_378_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_379_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_379_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_379_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_379_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_380_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_380_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_380_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_380_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_381_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_381_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_381_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_381_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_382_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_382_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_382_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_382_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_383_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_383_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_383_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_383_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_384_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_384_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_384_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_384_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_385_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_385_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_385_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_385_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_386_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_386_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_386_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_386_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_387_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_387_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_387_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_387_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_388_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_388_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_388_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_388_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_389_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_389_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_389_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_389_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_390_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_390_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_390_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_390_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_391_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_391_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_391_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_391_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_392_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_392_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_392_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_392_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_393_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_393_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_393_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_393_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_394_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_394_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_394_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_394_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_395_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_395_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_395_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_395_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_396_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_396_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_396_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_396_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_397_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_397_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_397_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_397_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_398_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_398_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_398_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_398_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_399_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_399_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_399_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_399_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_400_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_400_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_400_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_400_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_401_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_401_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_401_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_401_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_402_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_402_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_402_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_402_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_403_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_403_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_403_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_403_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_404_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_404_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_404_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_404_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_405_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_405_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_405_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_405_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_406_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_406_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_406_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_406_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_407_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_407_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_407_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_407_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_408_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_408_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_408_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_408_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_409_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_409_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_409_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_409_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_410_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_410_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_410_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_410_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_411_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_411_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_411_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_411_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_412_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_412_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_412_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_412_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_413_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_413_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_413_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_413_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_414_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_414_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_414_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_414_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_415_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_415_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_415_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_415_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_416_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_416_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_416_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_416_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_417_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_417_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_417_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_417_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_418_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_418_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_418_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_418_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_419_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_419_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_419_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_419_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_420_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_420_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_420_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_420_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_421_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_421_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_421_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_421_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_422_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_422_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_422_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_422_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_423_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_423_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_423_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_423_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_424_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_424_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_424_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_424_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_425_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_425_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_425_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_425_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_426_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_426_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_426_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_426_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_427_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_427_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_427_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_427_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_428_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_428_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_428_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_428_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_429_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_429_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_429_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_429_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_430_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_430_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_430_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_430_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_431_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_431_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_431_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_431_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_432_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_432_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_432_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_432_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_433_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_433_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_433_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_433_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_434_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_434_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_434_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_434_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_435_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_435_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_435_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_435_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_436_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_436_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_436_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_436_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_437_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_437_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_437_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_437_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_438_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_438_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_438_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_438_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_439_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_439_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_439_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_439_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_440_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_440_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_440_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_440_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_441_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_441_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_441_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_441_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_442_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_442_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_442_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_442_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_443_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_443_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_443_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_443_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_444_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_444_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_444_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_444_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_445_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_445_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_445_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_445_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_446_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_446_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_446_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_446_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_447_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_447_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_447_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_447_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_448_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_448_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_448_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_448_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_449_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_449_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_449_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_449_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_450_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_450_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_450_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_450_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_451_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_451_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_451_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_451_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_452_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_452_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_452_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_452_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_453_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_453_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_453_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_453_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_454_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_454_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_454_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_454_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_455_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_455_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_455_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_455_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_456_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_456_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_456_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_456_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_457_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_457_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_457_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_457_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_458_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_458_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_458_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_458_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_459_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_459_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_459_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_459_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_460_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_460_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_460_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_460_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_461_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_461_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_461_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_461_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_462_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_462_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_462_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_462_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_463_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_463_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_463_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_463_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_464_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_464_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_464_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_464_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_465_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_465_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_465_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_465_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_466_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_466_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_466_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_466_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_467_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_467_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_467_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_467_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_468_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_468_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_468_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_468_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_469_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_469_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_469_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_469_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_470_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_470_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_470_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_470_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_471_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_471_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_471_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_471_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_472_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_472_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_472_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_472_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_473_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_473_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_473_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_473_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_474_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_474_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_474_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_474_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_475_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_475_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_475_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_475_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_476_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_476_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_476_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_476_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_477_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_477_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_477_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_477_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_478_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_478_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_478_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_478_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_479_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_479_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_479_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_479_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_480_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_480_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_480_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_480_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_481_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_481_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_481_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_481_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_482_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_482_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_482_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_482_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_483_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_483_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_483_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_483_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_484_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_484_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_484_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_484_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_485_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_485_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_485_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_485_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_486_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_486_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_486_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_486_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_487_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_487_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_487_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_487_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_488_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_488_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_488_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_488_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_489_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_489_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_489_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_489_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_490_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_490_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_490_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_490_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_491_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_491_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_491_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_491_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_492_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_492_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_492_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_492_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_493_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_493_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_493_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_493_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_494_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_494_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_494_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_494_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_495_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_495_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_495_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_495_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_496_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_496_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_496_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_496_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_497_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_497_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_497_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_497_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_498_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_498_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_498_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_498_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_499_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_499_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_499_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_499_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_500_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_500_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_500_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_500_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_501_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_501_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_501_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_501_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_502_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_502_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_502_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_502_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_503_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_503_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_503_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_503_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_504_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_504_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_504_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_504_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_505_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_505_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_505_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_505_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_506_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_506_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_506_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_506_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_507_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_507_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_507_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_507_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_508_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_508_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_508_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_508_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_509_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_509_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_509_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_509_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_510_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_510_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_510_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_510_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_511_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_511_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_511_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_511_en; // @[SRAM_1.scala 63:26]
  wire [1:0] mem_MPORT_512_data; // @[SRAM_1.scala 63:26]
  wire [8:0] mem_MPORT_512_addr; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_512_mask; // @[SRAM_1.scala 63:26]
  wire  mem_MPORT_512_en; // @[SRAM_1.scala 63:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [8:0] mem_io_r_data_MPORT_addr_pipe_0;
  wire  readConflict = io_w_addr == io_r_addr; // @[SRAM_1.scala 81:34]
  assign mem_io_r_data_MPORT_en = mem_io_r_data_MPORT_en_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[SRAM_1.scala 63:26]
  assign mem_MPORT_data = 2'h0;
  assign mem_MPORT_addr = 9'h0;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = reset;
  assign mem_MPORT_1_data = 2'h0;
  assign mem_MPORT_1_addr = 9'h1;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = reset;
  assign mem_MPORT_2_data = 2'h0;
  assign mem_MPORT_2_addr = 9'h2;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = reset;
  assign mem_MPORT_3_data = 2'h0;
  assign mem_MPORT_3_addr = 9'h3;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = reset;
  assign mem_MPORT_4_data = 2'h0;
  assign mem_MPORT_4_addr = 9'h4;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = reset;
  assign mem_MPORT_5_data = 2'h0;
  assign mem_MPORT_5_addr = 9'h5;
  assign mem_MPORT_5_mask = 1'h1;
  assign mem_MPORT_5_en = reset;
  assign mem_MPORT_6_data = 2'h0;
  assign mem_MPORT_6_addr = 9'h6;
  assign mem_MPORT_6_mask = 1'h1;
  assign mem_MPORT_6_en = reset;
  assign mem_MPORT_7_data = 2'h0;
  assign mem_MPORT_7_addr = 9'h7;
  assign mem_MPORT_7_mask = 1'h1;
  assign mem_MPORT_7_en = reset;
  assign mem_MPORT_8_data = 2'h0;
  assign mem_MPORT_8_addr = 9'h8;
  assign mem_MPORT_8_mask = 1'h1;
  assign mem_MPORT_8_en = reset;
  assign mem_MPORT_9_data = 2'h0;
  assign mem_MPORT_9_addr = 9'h9;
  assign mem_MPORT_9_mask = 1'h1;
  assign mem_MPORT_9_en = reset;
  assign mem_MPORT_10_data = 2'h0;
  assign mem_MPORT_10_addr = 9'ha;
  assign mem_MPORT_10_mask = 1'h1;
  assign mem_MPORT_10_en = reset;
  assign mem_MPORT_11_data = 2'h0;
  assign mem_MPORT_11_addr = 9'hb;
  assign mem_MPORT_11_mask = 1'h1;
  assign mem_MPORT_11_en = reset;
  assign mem_MPORT_12_data = 2'h0;
  assign mem_MPORT_12_addr = 9'hc;
  assign mem_MPORT_12_mask = 1'h1;
  assign mem_MPORT_12_en = reset;
  assign mem_MPORT_13_data = 2'h0;
  assign mem_MPORT_13_addr = 9'hd;
  assign mem_MPORT_13_mask = 1'h1;
  assign mem_MPORT_13_en = reset;
  assign mem_MPORT_14_data = 2'h0;
  assign mem_MPORT_14_addr = 9'he;
  assign mem_MPORT_14_mask = 1'h1;
  assign mem_MPORT_14_en = reset;
  assign mem_MPORT_15_data = 2'h0;
  assign mem_MPORT_15_addr = 9'hf;
  assign mem_MPORT_15_mask = 1'h1;
  assign mem_MPORT_15_en = reset;
  assign mem_MPORT_16_data = 2'h0;
  assign mem_MPORT_16_addr = 9'h10;
  assign mem_MPORT_16_mask = 1'h1;
  assign mem_MPORT_16_en = reset;
  assign mem_MPORT_17_data = 2'h0;
  assign mem_MPORT_17_addr = 9'h11;
  assign mem_MPORT_17_mask = 1'h1;
  assign mem_MPORT_17_en = reset;
  assign mem_MPORT_18_data = 2'h0;
  assign mem_MPORT_18_addr = 9'h12;
  assign mem_MPORT_18_mask = 1'h1;
  assign mem_MPORT_18_en = reset;
  assign mem_MPORT_19_data = 2'h0;
  assign mem_MPORT_19_addr = 9'h13;
  assign mem_MPORT_19_mask = 1'h1;
  assign mem_MPORT_19_en = reset;
  assign mem_MPORT_20_data = 2'h0;
  assign mem_MPORT_20_addr = 9'h14;
  assign mem_MPORT_20_mask = 1'h1;
  assign mem_MPORT_20_en = reset;
  assign mem_MPORT_21_data = 2'h0;
  assign mem_MPORT_21_addr = 9'h15;
  assign mem_MPORT_21_mask = 1'h1;
  assign mem_MPORT_21_en = reset;
  assign mem_MPORT_22_data = 2'h0;
  assign mem_MPORT_22_addr = 9'h16;
  assign mem_MPORT_22_mask = 1'h1;
  assign mem_MPORT_22_en = reset;
  assign mem_MPORT_23_data = 2'h0;
  assign mem_MPORT_23_addr = 9'h17;
  assign mem_MPORT_23_mask = 1'h1;
  assign mem_MPORT_23_en = reset;
  assign mem_MPORT_24_data = 2'h0;
  assign mem_MPORT_24_addr = 9'h18;
  assign mem_MPORT_24_mask = 1'h1;
  assign mem_MPORT_24_en = reset;
  assign mem_MPORT_25_data = 2'h0;
  assign mem_MPORT_25_addr = 9'h19;
  assign mem_MPORT_25_mask = 1'h1;
  assign mem_MPORT_25_en = reset;
  assign mem_MPORT_26_data = 2'h0;
  assign mem_MPORT_26_addr = 9'h1a;
  assign mem_MPORT_26_mask = 1'h1;
  assign mem_MPORT_26_en = reset;
  assign mem_MPORT_27_data = 2'h0;
  assign mem_MPORT_27_addr = 9'h1b;
  assign mem_MPORT_27_mask = 1'h1;
  assign mem_MPORT_27_en = reset;
  assign mem_MPORT_28_data = 2'h0;
  assign mem_MPORT_28_addr = 9'h1c;
  assign mem_MPORT_28_mask = 1'h1;
  assign mem_MPORT_28_en = reset;
  assign mem_MPORT_29_data = 2'h0;
  assign mem_MPORT_29_addr = 9'h1d;
  assign mem_MPORT_29_mask = 1'h1;
  assign mem_MPORT_29_en = reset;
  assign mem_MPORT_30_data = 2'h0;
  assign mem_MPORT_30_addr = 9'h1e;
  assign mem_MPORT_30_mask = 1'h1;
  assign mem_MPORT_30_en = reset;
  assign mem_MPORT_31_data = 2'h0;
  assign mem_MPORT_31_addr = 9'h1f;
  assign mem_MPORT_31_mask = 1'h1;
  assign mem_MPORT_31_en = reset;
  assign mem_MPORT_32_data = 2'h0;
  assign mem_MPORT_32_addr = 9'h20;
  assign mem_MPORT_32_mask = 1'h1;
  assign mem_MPORT_32_en = reset;
  assign mem_MPORT_33_data = 2'h0;
  assign mem_MPORT_33_addr = 9'h21;
  assign mem_MPORT_33_mask = 1'h1;
  assign mem_MPORT_33_en = reset;
  assign mem_MPORT_34_data = 2'h0;
  assign mem_MPORT_34_addr = 9'h22;
  assign mem_MPORT_34_mask = 1'h1;
  assign mem_MPORT_34_en = reset;
  assign mem_MPORT_35_data = 2'h0;
  assign mem_MPORT_35_addr = 9'h23;
  assign mem_MPORT_35_mask = 1'h1;
  assign mem_MPORT_35_en = reset;
  assign mem_MPORT_36_data = 2'h0;
  assign mem_MPORT_36_addr = 9'h24;
  assign mem_MPORT_36_mask = 1'h1;
  assign mem_MPORT_36_en = reset;
  assign mem_MPORT_37_data = 2'h0;
  assign mem_MPORT_37_addr = 9'h25;
  assign mem_MPORT_37_mask = 1'h1;
  assign mem_MPORT_37_en = reset;
  assign mem_MPORT_38_data = 2'h0;
  assign mem_MPORT_38_addr = 9'h26;
  assign mem_MPORT_38_mask = 1'h1;
  assign mem_MPORT_38_en = reset;
  assign mem_MPORT_39_data = 2'h0;
  assign mem_MPORT_39_addr = 9'h27;
  assign mem_MPORT_39_mask = 1'h1;
  assign mem_MPORT_39_en = reset;
  assign mem_MPORT_40_data = 2'h0;
  assign mem_MPORT_40_addr = 9'h28;
  assign mem_MPORT_40_mask = 1'h1;
  assign mem_MPORT_40_en = reset;
  assign mem_MPORT_41_data = 2'h0;
  assign mem_MPORT_41_addr = 9'h29;
  assign mem_MPORT_41_mask = 1'h1;
  assign mem_MPORT_41_en = reset;
  assign mem_MPORT_42_data = 2'h0;
  assign mem_MPORT_42_addr = 9'h2a;
  assign mem_MPORT_42_mask = 1'h1;
  assign mem_MPORT_42_en = reset;
  assign mem_MPORT_43_data = 2'h0;
  assign mem_MPORT_43_addr = 9'h2b;
  assign mem_MPORT_43_mask = 1'h1;
  assign mem_MPORT_43_en = reset;
  assign mem_MPORT_44_data = 2'h0;
  assign mem_MPORT_44_addr = 9'h2c;
  assign mem_MPORT_44_mask = 1'h1;
  assign mem_MPORT_44_en = reset;
  assign mem_MPORT_45_data = 2'h0;
  assign mem_MPORT_45_addr = 9'h2d;
  assign mem_MPORT_45_mask = 1'h1;
  assign mem_MPORT_45_en = reset;
  assign mem_MPORT_46_data = 2'h0;
  assign mem_MPORT_46_addr = 9'h2e;
  assign mem_MPORT_46_mask = 1'h1;
  assign mem_MPORT_46_en = reset;
  assign mem_MPORT_47_data = 2'h0;
  assign mem_MPORT_47_addr = 9'h2f;
  assign mem_MPORT_47_mask = 1'h1;
  assign mem_MPORT_47_en = reset;
  assign mem_MPORT_48_data = 2'h0;
  assign mem_MPORT_48_addr = 9'h30;
  assign mem_MPORT_48_mask = 1'h1;
  assign mem_MPORT_48_en = reset;
  assign mem_MPORT_49_data = 2'h0;
  assign mem_MPORT_49_addr = 9'h31;
  assign mem_MPORT_49_mask = 1'h1;
  assign mem_MPORT_49_en = reset;
  assign mem_MPORT_50_data = 2'h0;
  assign mem_MPORT_50_addr = 9'h32;
  assign mem_MPORT_50_mask = 1'h1;
  assign mem_MPORT_50_en = reset;
  assign mem_MPORT_51_data = 2'h0;
  assign mem_MPORT_51_addr = 9'h33;
  assign mem_MPORT_51_mask = 1'h1;
  assign mem_MPORT_51_en = reset;
  assign mem_MPORT_52_data = 2'h0;
  assign mem_MPORT_52_addr = 9'h34;
  assign mem_MPORT_52_mask = 1'h1;
  assign mem_MPORT_52_en = reset;
  assign mem_MPORT_53_data = 2'h0;
  assign mem_MPORT_53_addr = 9'h35;
  assign mem_MPORT_53_mask = 1'h1;
  assign mem_MPORT_53_en = reset;
  assign mem_MPORT_54_data = 2'h0;
  assign mem_MPORT_54_addr = 9'h36;
  assign mem_MPORT_54_mask = 1'h1;
  assign mem_MPORT_54_en = reset;
  assign mem_MPORT_55_data = 2'h0;
  assign mem_MPORT_55_addr = 9'h37;
  assign mem_MPORT_55_mask = 1'h1;
  assign mem_MPORT_55_en = reset;
  assign mem_MPORT_56_data = 2'h0;
  assign mem_MPORT_56_addr = 9'h38;
  assign mem_MPORT_56_mask = 1'h1;
  assign mem_MPORT_56_en = reset;
  assign mem_MPORT_57_data = 2'h0;
  assign mem_MPORT_57_addr = 9'h39;
  assign mem_MPORT_57_mask = 1'h1;
  assign mem_MPORT_57_en = reset;
  assign mem_MPORT_58_data = 2'h0;
  assign mem_MPORT_58_addr = 9'h3a;
  assign mem_MPORT_58_mask = 1'h1;
  assign mem_MPORT_58_en = reset;
  assign mem_MPORT_59_data = 2'h0;
  assign mem_MPORT_59_addr = 9'h3b;
  assign mem_MPORT_59_mask = 1'h1;
  assign mem_MPORT_59_en = reset;
  assign mem_MPORT_60_data = 2'h0;
  assign mem_MPORT_60_addr = 9'h3c;
  assign mem_MPORT_60_mask = 1'h1;
  assign mem_MPORT_60_en = reset;
  assign mem_MPORT_61_data = 2'h0;
  assign mem_MPORT_61_addr = 9'h3d;
  assign mem_MPORT_61_mask = 1'h1;
  assign mem_MPORT_61_en = reset;
  assign mem_MPORT_62_data = 2'h0;
  assign mem_MPORT_62_addr = 9'h3e;
  assign mem_MPORT_62_mask = 1'h1;
  assign mem_MPORT_62_en = reset;
  assign mem_MPORT_63_data = 2'h0;
  assign mem_MPORT_63_addr = 9'h3f;
  assign mem_MPORT_63_mask = 1'h1;
  assign mem_MPORT_63_en = reset;
  assign mem_MPORT_64_data = 2'h0;
  assign mem_MPORT_64_addr = 9'h40;
  assign mem_MPORT_64_mask = 1'h1;
  assign mem_MPORT_64_en = reset;
  assign mem_MPORT_65_data = 2'h0;
  assign mem_MPORT_65_addr = 9'h41;
  assign mem_MPORT_65_mask = 1'h1;
  assign mem_MPORT_65_en = reset;
  assign mem_MPORT_66_data = 2'h0;
  assign mem_MPORT_66_addr = 9'h42;
  assign mem_MPORT_66_mask = 1'h1;
  assign mem_MPORT_66_en = reset;
  assign mem_MPORT_67_data = 2'h0;
  assign mem_MPORT_67_addr = 9'h43;
  assign mem_MPORT_67_mask = 1'h1;
  assign mem_MPORT_67_en = reset;
  assign mem_MPORT_68_data = 2'h0;
  assign mem_MPORT_68_addr = 9'h44;
  assign mem_MPORT_68_mask = 1'h1;
  assign mem_MPORT_68_en = reset;
  assign mem_MPORT_69_data = 2'h0;
  assign mem_MPORT_69_addr = 9'h45;
  assign mem_MPORT_69_mask = 1'h1;
  assign mem_MPORT_69_en = reset;
  assign mem_MPORT_70_data = 2'h0;
  assign mem_MPORT_70_addr = 9'h46;
  assign mem_MPORT_70_mask = 1'h1;
  assign mem_MPORT_70_en = reset;
  assign mem_MPORT_71_data = 2'h0;
  assign mem_MPORT_71_addr = 9'h47;
  assign mem_MPORT_71_mask = 1'h1;
  assign mem_MPORT_71_en = reset;
  assign mem_MPORT_72_data = 2'h0;
  assign mem_MPORT_72_addr = 9'h48;
  assign mem_MPORT_72_mask = 1'h1;
  assign mem_MPORT_72_en = reset;
  assign mem_MPORT_73_data = 2'h0;
  assign mem_MPORT_73_addr = 9'h49;
  assign mem_MPORT_73_mask = 1'h1;
  assign mem_MPORT_73_en = reset;
  assign mem_MPORT_74_data = 2'h0;
  assign mem_MPORT_74_addr = 9'h4a;
  assign mem_MPORT_74_mask = 1'h1;
  assign mem_MPORT_74_en = reset;
  assign mem_MPORT_75_data = 2'h0;
  assign mem_MPORT_75_addr = 9'h4b;
  assign mem_MPORT_75_mask = 1'h1;
  assign mem_MPORT_75_en = reset;
  assign mem_MPORT_76_data = 2'h0;
  assign mem_MPORT_76_addr = 9'h4c;
  assign mem_MPORT_76_mask = 1'h1;
  assign mem_MPORT_76_en = reset;
  assign mem_MPORT_77_data = 2'h0;
  assign mem_MPORT_77_addr = 9'h4d;
  assign mem_MPORT_77_mask = 1'h1;
  assign mem_MPORT_77_en = reset;
  assign mem_MPORT_78_data = 2'h0;
  assign mem_MPORT_78_addr = 9'h4e;
  assign mem_MPORT_78_mask = 1'h1;
  assign mem_MPORT_78_en = reset;
  assign mem_MPORT_79_data = 2'h0;
  assign mem_MPORT_79_addr = 9'h4f;
  assign mem_MPORT_79_mask = 1'h1;
  assign mem_MPORT_79_en = reset;
  assign mem_MPORT_80_data = 2'h0;
  assign mem_MPORT_80_addr = 9'h50;
  assign mem_MPORT_80_mask = 1'h1;
  assign mem_MPORT_80_en = reset;
  assign mem_MPORT_81_data = 2'h0;
  assign mem_MPORT_81_addr = 9'h51;
  assign mem_MPORT_81_mask = 1'h1;
  assign mem_MPORT_81_en = reset;
  assign mem_MPORT_82_data = 2'h0;
  assign mem_MPORT_82_addr = 9'h52;
  assign mem_MPORT_82_mask = 1'h1;
  assign mem_MPORT_82_en = reset;
  assign mem_MPORT_83_data = 2'h0;
  assign mem_MPORT_83_addr = 9'h53;
  assign mem_MPORT_83_mask = 1'h1;
  assign mem_MPORT_83_en = reset;
  assign mem_MPORT_84_data = 2'h0;
  assign mem_MPORT_84_addr = 9'h54;
  assign mem_MPORT_84_mask = 1'h1;
  assign mem_MPORT_84_en = reset;
  assign mem_MPORT_85_data = 2'h0;
  assign mem_MPORT_85_addr = 9'h55;
  assign mem_MPORT_85_mask = 1'h1;
  assign mem_MPORT_85_en = reset;
  assign mem_MPORT_86_data = 2'h0;
  assign mem_MPORT_86_addr = 9'h56;
  assign mem_MPORT_86_mask = 1'h1;
  assign mem_MPORT_86_en = reset;
  assign mem_MPORT_87_data = 2'h0;
  assign mem_MPORT_87_addr = 9'h57;
  assign mem_MPORT_87_mask = 1'h1;
  assign mem_MPORT_87_en = reset;
  assign mem_MPORT_88_data = 2'h0;
  assign mem_MPORT_88_addr = 9'h58;
  assign mem_MPORT_88_mask = 1'h1;
  assign mem_MPORT_88_en = reset;
  assign mem_MPORT_89_data = 2'h0;
  assign mem_MPORT_89_addr = 9'h59;
  assign mem_MPORT_89_mask = 1'h1;
  assign mem_MPORT_89_en = reset;
  assign mem_MPORT_90_data = 2'h0;
  assign mem_MPORT_90_addr = 9'h5a;
  assign mem_MPORT_90_mask = 1'h1;
  assign mem_MPORT_90_en = reset;
  assign mem_MPORT_91_data = 2'h0;
  assign mem_MPORT_91_addr = 9'h5b;
  assign mem_MPORT_91_mask = 1'h1;
  assign mem_MPORT_91_en = reset;
  assign mem_MPORT_92_data = 2'h0;
  assign mem_MPORT_92_addr = 9'h5c;
  assign mem_MPORT_92_mask = 1'h1;
  assign mem_MPORT_92_en = reset;
  assign mem_MPORT_93_data = 2'h0;
  assign mem_MPORT_93_addr = 9'h5d;
  assign mem_MPORT_93_mask = 1'h1;
  assign mem_MPORT_93_en = reset;
  assign mem_MPORT_94_data = 2'h0;
  assign mem_MPORT_94_addr = 9'h5e;
  assign mem_MPORT_94_mask = 1'h1;
  assign mem_MPORT_94_en = reset;
  assign mem_MPORT_95_data = 2'h0;
  assign mem_MPORT_95_addr = 9'h5f;
  assign mem_MPORT_95_mask = 1'h1;
  assign mem_MPORT_95_en = reset;
  assign mem_MPORT_96_data = 2'h0;
  assign mem_MPORT_96_addr = 9'h60;
  assign mem_MPORT_96_mask = 1'h1;
  assign mem_MPORT_96_en = reset;
  assign mem_MPORT_97_data = 2'h0;
  assign mem_MPORT_97_addr = 9'h61;
  assign mem_MPORT_97_mask = 1'h1;
  assign mem_MPORT_97_en = reset;
  assign mem_MPORT_98_data = 2'h0;
  assign mem_MPORT_98_addr = 9'h62;
  assign mem_MPORT_98_mask = 1'h1;
  assign mem_MPORT_98_en = reset;
  assign mem_MPORT_99_data = 2'h0;
  assign mem_MPORT_99_addr = 9'h63;
  assign mem_MPORT_99_mask = 1'h1;
  assign mem_MPORT_99_en = reset;
  assign mem_MPORT_100_data = 2'h0;
  assign mem_MPORT_100_addr = 9'h64;
  assign mem_MPORT_100_mask = 1'h1;
  assign mem_MPORT_100_en = reset;
  assign mem_MPORT_101_data = 2'h0;
  assign mem_MPORT_101_addr = 9'h65;
  assign mem_MPORT_101_mask = 1'h1;
  assign mem_MPORT_101_en = reset;
  assign mem_MPORT_102_data = 2'h0;
  assign mem_MPORT_102_addr = 9'h66;
  assign mem_MPORT_102_mask = 1'h1;
  assign mem_MPORT_102_en = reset;
  assign mem_MPORT_103_data = 2'h0;
  assign mem_MPORT_103_addr = 9'h67;
  assign mem_MPORT_103_mask = 1'h1;
  assign mem_MPORT_103_en = reset;
  assign mem_MPORT_104_data = 2'h0;
  assign mem_MPORT_104_addr = 9'h68;
  assign mem_MPORT_104_mask = 1'h1;
  assign mem_MPORT_104_en = reset;
  assign mem_MPORT_105_data = 2'h0;
  assign mem_MPORT_105_addr = 9'h69;
  assign mem_MPORT_105_mask = 1'h1;
  assign mem_MPORT_105_en = reset;
  assign mem_MPORT_106_data = 2'h0;
  assign mem_MPORT_106_addr = 9'h6a;
  assign mem_MPORT_106_mask = 1'h1;
  assign mem_MPORT_106_en = reset;
  assign mem_MPORT_107_data = 2'h0;
  assign mem_MPORT_107_addr = 9'h6b;
  assign mem_MPORT_107_mask = 1'h1;
  assign mem_MPORT_107_en = reset;
  assign mem_MPORT_108_data = 2'h0;
  assign mem_MPORT_108_addr = 9'h6c;
  assign mem_MPORT_108_mask = 1'h1;
  assign mem_MPORT_108_en = reset;
  assign mem_MPORT_109_data = 2'h0;
  assign mem_MPORT_109_addr = 9'h6d;
  assign mem_MPORT_109_mask = 1'h1;
  assign mem_MPORT_109_en = reset;
  assign mem_MPORT_110_data = 2'h0;
  assign mem_MPORT_110_addr = 9'h6e;
  assign mem_MPORT_110_mask = 1'h1;
  assign mem_MPORT_110_en = reset;
  assign mem_MPORT_111_data = 2'h0;
  assign mem_MPORT_111_addr = 9'h6f;
  assign mem_MPORT_111_mask = 1'h1;
  assign mem_MPORT_111_en = reset;
  assign mem_MPORT_112_data = 2'h0;
  assign mem_MPORT_112_addr = 9'h70;
  assign mem_MPORT_112_mask = 1'h1;
  assign mem_MPORT_112_en = reset;
  assign mem_MPORT_113_data = 2'h0;
  assign mem_MPORT_113_addr = 9'h71;
  assign mem_MPORT_113_mask = 1'h1;
  assign mem_MPORT_113_en = reset;
  assign mem_MPORT_114_data = 2'h0;
  assign mem_MPORT_114_addr = 9'h72;
  assign mem_MPORT_114_mask = 1'h1;
  assign mem_MPORT_114_en = reset;
  assign mem_MPORT_115_data = 2'h0;
  assign mem_MPORT_115_addr = 9'h73;
  assign mem_MPORT_115_mask = 1'h1;
  assign mem_MPORT_115_en = reset;
  assign mem_MPORT_116_data = 2'h0;
  assign mem_MPORT_116_addr = 9'h74;
  assign mem_MPORT_116_mask = 1'h1;
  assign mem_MPORT_116_en = reset;
  assign mem_MPORT_117_data = 2'h0;
  assign mem_MPORT_117_addr = 9'h75;
  assign mem_MPORT_117_mask = 1'h1;
  assign mem_MPORT_117_en = reset;
  assign mem_MPORT_118_data = 2'h0;
  assign mem_MPORT_118_addr = 9'h76;
  assign mem_MPORT_118_mask = 1'h1;
  assign mem_MPORT_118_en = reset;
  assign mem_MPORT_119_data = 2'h0;
  assign mem_MPORT_119_addr = 9'h77;
  assign mem_MPORT_119_mask = 1'h1;
  assign mem_MPORT_119_en = reset;
  assign mem_MPORT_120_data = 2'h0;
  assign mem_MPORT_120_addr = 9'h78;
  assign mem_MPORT_120_mask = 1'h1;
  assign mem_MPORT_120_en = reset;
  assign mem_MPORT_121_data = 2'h0;
  assign mem_MPORT_121_addr = 9'h79;
  assign mem_MPORT_121_mask = 1'h1;
  assign mem_MPORT_121_en = reset;
  assign mem_MPORT_122_data = 2'h0;
  assign mem_MPORT_122_addr = 9'h7a;
  assign mem_MPORT_122_mask = 1'h1;
  assign mem_MPORT_122_en = reset;
  assign mem_MPORT_123_data = 2'h0;
  assign mem_MPORT_123_addr = 9'h7b;
  assign mem_MPORT_123_mask = 1'h1;
  assign mem_MPORT_123_en = reset;
  assign mem_MPORT_124_data = 2'h0;
  assign mem_MPORT_124_addr = 9'h7c;
  assign mem_MPORT_124_mask = 1'h1;
  assign mem_MPORT_124_en = reset;
  assign mem_MPORT_125_data = 2'h0;
  assign mem_MPORT_125_addr = 9'h7d;
  assign mem_MPORT_125_mask = 1'h1;
  assign mem_MPORT_125_en = reset;
  assign mem_MPORT_126_data = 2'h0;
  assign mem_MPORT_126_addr = 9'h7e;
  assign mem_MPORT_126_mask = 1'h1;
  assign mem_MPORT_126_en = reset;
  assign mem_MPORT_127_data = 2'h0;
  assign mem_MPORT_127_addr = 9'h7f;
  assign mem_MPORT_127_mask = 1'h1;
  assign mem_MPORT_127_en = reset;
  assign mem_MPORT_128_data = 2'h0;
  assign mem_MPORT_128_addr = 9'h80;
  assign mem_MPORT_128_mask = 1'h1;
  assign mem_MPORT_128_en = reset;
  assign mem_MPORT_129_data = 2'h0;
  assign mem_MPORT_129_addr = 9'h81;
  assign mem_MPORT_129_mask = 1'h1;
  assign mem_MPORT_129_en = reset;
  assign mem_MPORT_130_data = 2'h0;
  assign mem_MPORT_130_addr = 9'h82;
  assign mem_MPORT_130_mask = 1'h1;
  assign mem_MPORT_130_en = reset;
  assign mem_MPORT_131_data = 2'h0;
  assign mem_MPORT_131_addr = 9'h83;
  assign mem_MPORT_131_mask = 1'h1;
  assign mem_MPORT_131_en = reset;
  assign mem_MPORT_132_data = 2'h0;
  assign mem_MPORT_132_addr = 9'h84;
  assign mem_MPORT_132_mask = 1'h1;
  assign mem_MPORT_132_en = reset;
  assign mem_MPORT_133_data = 2'h0;
  assign mem_MPORT_133_addr = 9'h85;
  assign mem_MPORT_133_mask = 1'h1;
  assign mem_MPORT_133_en = reset;
  assign mem_MPORT_134_data = 2'h0;
  assign mem_MPORT_134_addr = 9'h86;
  assign mem_MPORT_134_mask = 1'h1;
  assign mem_MPORT_134_en = reset;
  assign mem_MPORT_135_data = 2'h0;
  assign mem_MPORT_135_addr = 9'h87;
  assign mem_MPORT_135_mask = 1'h1;
  assign mem_MPORT_135_en = reset;
  assign mem_MPORT_136_data = 2'h0;
  assign mem_MPORT_136_addr = 9'h88;
  assign mem_MPORT_136_mask = 1'h1;
  assign mem_MPORT_136_en = reset;
  assign mem_MPORT_137_data = 2'h0;
  assign mem_MPORT_137_addr = 9'h89;
  assign mem_MPORT_137_mask = 1'h1;
  assign mem_MPORT_137_en = reset;
  assign mem_MPORT_138_data = 2'h0;
  assign mem_MPORT_138_addr = 9'h8a;
  assign mem_MPORT_138_mask = 1'h1;
  assign mem_MPORT_138_en = reset;
  assign mem_MPORT_139_data = 2'h0;
  assign mem_MPORT_139_addr = 9'h8b;
  assign mem_MPORT_139_mask = 1'h1;
  assign mem_MPORT_139_en = reset;
  assign mem_MPORT_140_data = 2'h0;
  assign mem_MPORT_140_addr = 9'h8c;
  assign mem_MPORT_140_mask = 1'h1;
  assign mem_MPORT_140_en = reset;
  assign mem_MPORT_141_data = 2'h0;
  assign mem_MPORT_141_addr = 9'h8d;
  assign mem_MPORT_141_mask = 1'h1;
  assign mem_MPORT_141_en = reset;
  assign mem_MPORT_142_data = 2'h0;
  assign mem_MPORT_142_addr = 9'h8e;
  assign mem_MPORT_142_mask = 1'h1;
  assign mem_MPORT_142_en = reset;
  assign mem_MPORT_143_data = 2'h0;
  assign mem_MPORT_143_addr = 9'h8f;
  assign mem_MPORT_143_mask = 1'h1;
  assign mem_MPORT_143_en = reset;
  assign mem_MPORT_144_data = 2'h0;
  assign mem_MPORT_144_addr = 9'h90;
  assign mem_MPORT_144_mask = 1'h1;
  assign mem_MPORT_144_en = reset;
  assign mem_MPORT_145_data = 2'h0;
  assign mem_MPORT_145_addr = 9'h91;
  assign mem_MPORT_145_mask = 1'h1;
  assign mem_MPORT_145_en = reset;
  assign mem_MPORT_146_data = 2'h0;
  assign mem_MPORT_146_addr = 9'h92;
  assign mem_MPORT_146_mask = 1'h1;
  assign mem_MPORT_146_en = reset;
  assign mem_MPORT_147_data = 2'h0;
  assign mem_MPORT_147_addr = 9'h93;
  assign mem_MPORT_147_mask = 1'h1;
  assign mem_MPORT_147_en = reset;
  assign mem_MPORT_148_data = 2'h0;
  assign mem_MPORT_148_addr = 9'h94;
  assign mem_MPORT_148_mask = 1'h1;
  assign mem_MPORT_148_en = reset;
  assign mem_MPORT_149_data = 2'h0;
  assign mem_MPORT_149_addr = 9'h95;
  assign mem_MPORT_149_mask = 1'h1;
  assign mem_MPORT_149_en = reset;
  assign mem_MPORT_150_data = 2'h0;
  assign mem_MPORT_150_addr = 9'h96;
  assign mem_MPORT_150_mask = 1'h1;
  assign mem_MPORT_150_en = reset;
  assign mem_MPORT_151_data = 2'h0;
  assign mem_MPORT_151_addr = 9'h97;
  assign mem_MPORT_151_mask = 1'h1;
  assign mem_MPORT_151_en = reset;
  assign mem_MPORT_152_data = 2'h0;
  assign mem_MPORT_152_addr = 9'h98;
  assign mem_MPORT_152_mask = 1'h1;
  assign mem_MPORT_152_en = reset;
  assign mem_MPORT_153_data = 2'h0;
  assign mem_MPORT_153_addr = 9'h99;
  assign mem_MPORT_153_mask = 1'h1;
  assign mem_MPORT_153_en = reset;
  assign mem_MPORT_154_data = 2'h0;
  assign mem_MPORT_154_addr = 9'h9a;
  assign mem_MPORT_154_mask = 1'h1;
  assign mem_MPORT_154_en = reset;
  assign mem_MPORT_155_data = 2'h0;
  assign mem_MPORT_155_addr = 9'h9b;
  assign mem_MPORT_155_mask = 1'h1;
  assign mem_MPORT_155_en = reset;
  assign mem_MPORT_156_data = 2'h0;
  assign mem_MPORT_156_addr = 9'h9c;
  assign mem_MPORT_156_mask = 1'h1;
  assign mem_MPORT_156_en = reset;
  assign mem_MPORT_157_data = 2'h0;
  assign mem_MPORT_157_addr = 9'h9d;
  assign mem_MPORT_157_mask = 1'h1;
  assign mem_MPORT_157_en = reset;
  assign mem_MPORT_158_data = 2'h0;
  assign mem_MPORT_158_addr = 9'h9e;
  assign mem_MPORT_158_mask = 1'h1;
  assign mem_MPORT_158_en = reset;
  assign mem_MPORT_159_data = 2'h0;
  assign mem_MPORT_159_addr = 9'h9f;
  assign mem_MPORT_159_mask = 1'h1;
  assign mem_MPORT_159_en = reset;
  assign mem_MPORT_160_data = 2'h0;
  assign mem_MPORT_160_addr = 9'ha0;
  assign mem_MPORT_160_mask = 1'h1;
  assign mem_MPORT_160_en = reset;
  assign mem_MPORT_161_data = 2'h0;
  assign mem_MPORT_161_addr = 9'ha1;
  assign mem_MPORT_161_mask = 1'h1;
  assign mem_MPORT_161_en = reset;
  assign mem_MPORT_162_data = 2'h0;
  assign mem_MPORT_162_addr = 9'ha2;
  assign mem_MPORT_162_mask = 1'h1;
  assign mem_MPORT_162_en = reset;
  assign mem_MPORT_163_data = 2'h0;
  assign mem_MPORT_163_addr = 9'ha3;
  assign mem_MPORT_163_mask = 1'h1;
  assign mem_MPORT_163_en = reset;
  assign mem_MPORT_164_data = 2'h0;
  assign mem_MPORT_164_addr = 9'ha4;
  assign mem_MPORT_164_mask = 1'h1;
  assign mem_MPORT_164_en = reset;
  assign mem_MPORT_165_data = 2'h0;
  assign mem_MPORT_165_addr = 9'ha5;
  assign mem_MPORT_165_mask = 1'h1;
  assign mem_MPORT_165_en = reset;
  assign mem_MPORT_166_data = 2'h0;
  assign mem_MPORT_166_addr = 9'ha6;
  assign mem_MPORT_166_mask = 1'h1;
  assign mem_MPORT_166_en = reset;
  assign mem_MPORT_167_data = 2'h0;
  assign mem_MPORT_167_addr = 9'ha7;
  assign mem_MPORT_167_mask = 1'h1;
  assign mem_MPORT_167_en = reset;
  assign mem_MPORT_168_data = 2'h0;
  assign mem_MPORT_168_addr = 9'ha8;
  assign mem_MPORT_168_mask = 1'h1;
  assign mem_MPORT_168_en = reset;
  assign mem_MPORT_169_data = 2'h0;
  assign mem_MPORT_169_addr = 9'ha9;
  assign mem_MPORT_169_mask = 1'h1;
  assign mem_MPORT_169_en = reset;
  assign mem_MPORT_170_data = 2'h0;
  assign mem_MPORT_170_addr = 9'haa;
  assign mem_MPORT_170_mask = 1'h1;
  assign mem_MPORT_170_en = reset;
  assign mem_MPORT_171_data = 2'h0;
  assign mem_MPORT_171_addr = 9'hab;
  assign mem_MPORT_171_mask = 1'h1;
  assign mem_MPORT_171_en = reset;
  assign mem_MPORT_172_data = 2'h0;
  assign mem_MPORT_172_addr = 9'hac;
  assign mem_MPORT_172_mask = 1'h1;
  assign mem_MPORT_172_en = reset;
  assign mem_MPORT_173_data = 2'h0;
  assign mem_MPORT_173_addr = 9'had;
  assign mem_MPORT_173_mask = 1'h1;
  assign mem_MPORT_173_en = reset;
  assign mem_MPORT_174_data = 2'h0;
  assign mem_MPORT_174_addr = 9'hae;
  assign mem_MPORT_174_mask = 1'h1;
  assign mem_MPORT_174_en = reset;
  assign mem_MPORT_175_data = 2'h0;
  assign mem_MPORT_175_addr = 9'haf;
  assign mem_MPORT_175_mask = 1'h1;
  assign mem_MPORT_175_en = reset;
  assign mem_MPORT_176_data = 2'h0;
  assign mem_MPORT_176_addr = 9'hb0;
  assign mem_MPORT_176_mask = 1'h1;
  assign mem_MPORT_176_en = reset;
  assign mem_MPORT_177_data = 2'h0;
  assign mem_MPORT_177_addr = 9'hb1;
  assign mem_MPORT_177_mask = 1'h1;
  assign mem_MPORT_177_en = reset;
  assign mem_MPORT_178_data = 2'h0;
  assign mem_MPORT_178_addr = 9'hb2;
  assign mem_MPORT_178_mask = 1'h1;
  assign mem_MPORT_178_en = reset;
  assign mem_MPORT_179_data = 2'h0;
  assign mem_MPORT_179_addr = 9'hb3;
  assign mem_MPORT_179_mask = 1'h1;
  assign mem_MPORT_179_en = reset;
  assign mem_MPORT_180_data = 2'h0;
  assign mem_MPORT_180_addr = 9'hb4;
  assign mem_MPORT_180_mask = 1'h1;
  assign mem_MPORT_180_en = reset;
  assign mem_MPORT_181_data = 2'h0;
  assign mem_MPORT_181_addr = 9'hb5;
  assign mem_MPORT_181_mask = 1'h1;
  assign mem_MPORT_181_en = reset;
  assign mem_MPORT_182_data = 2'h0;
  assign mem_MPORT_182_addr = 9'hb6;
  assign mem_MPORT_182_mask = 1'h1;
  assign mem_MPORT_182_en = reset;
  assign mem_MPORT_183_data = 2'h0;
  assign mem_MPORT_183_addr = 9'hb7;
  assign mem_MPORT_183_mask = 1'h1;
  assign mem_MPORT_183_en = reset;
  assign mem_MPORT_184_data = 2'h0;
  assign mem_MPORT_184_addr = 9'hb8;
  assign mem_MPORT_184_mask = 1'h1;
  assign mem_MPORT_184_en = reset;
  assign mem_MPORT_185_data = 2'h0;
  assign mem_MPORT_185_addr = 9'hb9;
  assign mem_MPORT_185_mask = 1'h1;
  assign mem_MPORT_185_en = reset;
  assign mem_MPORT_186_data = 2'h0;
  assign mem_MPORT_186_addr = 9'hba;
  assign mem_MPORT_186_mask = 1'h1;
  assign mem_MPORT_186_en = reset;
  assign mem_MPORT_187_data = 2'h0;
  assign mem_MPORT_187_addr = 9'hbb;
  assign mem_MPORT_187_mask = 1'h1;
  assign mem_MPORT_187_en = reset;
  assign mem_MPORT_188_data = 2'h0;
  assign mem_MPORT_188_addr = 9'hbc;
  assign mem_MPORT_188_mask = 1'h1;
  assign mem_MPORT_188_en = reset;
  assign mem_MPORT_189_data = 2'h0;
  assign mem_MPORT_189_addr = 9'hbd;
  assign mem_MPORT_189_mask = 1'h1;
  assign mem_MPORT_189_en = reset;
  assign mem_MPORT_190_data = 2'h0;
  assign mem_MPORT_190_addr = 9'hbe;
  assign mem_MPORT_190_mask = 1'h1;
  assign mem_MPORT_190_en = reset;
  assign mem_MPORT_191_data = 2'h0;
  assign mem_MPORT_191_addr = 9'hbf;
  assign mem_MPORT_191_mask = 1'h1;
  assign mem_MPORT_191_en = reset;
  assign mem_MPORT_192_data = 2'h0;
  assign mem_MPORT_192_addr = 9'hc0;
  assign mem_MPORT_192_mask = 1'h1;
  assign mem_MPORT_192_en = reset;
  assign mem_MPORT_193_data = 2'h0;
  assign mem_MPORT_193_addr = 9'hc1;
  assign mem_MPORT_193_mask = 1'h1;
  assign mem_MPORT_193_en = reset;
  assign mem_MPORT_194_data = 2'h0;
  assign mem_MPORT_194_addr = 9'hc2;
  assign mem_MPORT_194_mask = 1'h1;
  assign mem_MPORT_194_en = reset;
  assign mem_MPORT_195_data = 2'h0;
  assign mem_MPORT_195_addr = 9'hc3;
  assign mem_MPORT_195_mask = 1'h1;
  assign mem_MPORT_195_en = reset;
  assign mem_MPORT_196_data = 2'h0;
  assign mem_MPORT_196_addr = 9'hc4;
  assign mem_MPORT_196_mask = 1'h1;
  assign mem_MPORT_196_en = reset;
  assign mem_MPORT_197_data = 2'h0;
  assign mem_MPORT_197_addr = 9'hc5;
  assign mem_MPORT_197_mask = 1'h1;
  assign mem_MPORT_197_en = reset;
  assign mem_MPORT_198_data = 2'h0;
  assign mem_MPORT_198_addr = 9'hc6;
  assign mem_MPORT_198_mask = 1'h1;
  assign mem_MPORT_198_en = reset;
  assign mem_MPORT_199_data = 2'h0;
  assign mem_MPORT_199_addr = 9'hc7;
  assign mem_MPORT_199_mask = 1'h1;
  assign mem_MPORT_199_en = reset;
  assign mem_MPORT_200_data = 2'h0;
  assign mem_MPORT_200_addr = 9'hc8;
  assign mem_MPORT_200_mask = 1'h1;
  assign mem_MPORT_200_en = reset;
  assign mem_MPORT_201_data = 2'h0;
  assign mem_MPORT_201_addr = 9'hc9;
  assign mem_MPORT_201_mask = 1'h1;
  assign mem_MPORT_201_en = reset;
  assign mem_MPORT_202_data = 2'h0;
  assign mem_MPORT_202_addr = 9'hca;
  assign mem_MPORT_202_mask = 1'h1;
  assign mem_MPORT_202_en = reset;
  assign mem_MPORT_203_data = 2'h0;
  assign mem_MPORT_203_addr = 9'hcb;
  assign mem_MPORT_203_mask = 1'h1;
  assign mem_MPORT_203_en = reset;
  assign mem_MPORT_204_data = 2'h0;
  assign mem_MPORT_204_addr = 9'hcc;
  assign mem_MPORT_204_mask = 1'h1;
  assign mem_MPORT_204_en = reset;
  assign mem_MPORT_205_data = 2'h0;
  assign mem_MPORT_205_addr = 9'hcd;
  assign mem_MPORT_205_mask = 1'h1;
  assign mem_MPORT_205_en = reset;
  assign mem_MPORT_206_data = 2'h0;
  assign mem_MPORT_206_addr = 9'hce;
  assign mem_MPORT_206_mask = 1'h1;
  assign mem_MPORT_206_en = reset;
  assign mem_MPORT_207_data = 2'h0;
  assign mem_MPORT_207_addr = 9'hcf;
  assign mem_MPORT_207_mask = 1'h1;
  assign mem_MPORT_207_en = reset;
  assign mem_MPORT_208_data = 2'h0;
  assign mem_MPORT_208_addr = 9'hd0;
  assign mem_MPORT_208_mask = 1'h1;
  assign mem_MPORT_208_en = reset;
  assign mem_MPORT_209_data = 2'h0;
  assign mem_MPORT_209_addr = 9'hd1;
  assign mem_MPORT_209_mask = 1'h1;
  assign mem_MPORT_209_en = reset;
  assign mem_MPORT_210_data = 2'h0;
  assign mem_MPORT_210_addr = 9'hd2;
  assign mem_MPORT_210_mask = 1'h1;
  assign mem_MPORT_210_en = reset;
  assign mem_MPORT_211_data = 2'h0;
  assign mem_MPORT_211_addr = 9'hd3;
  assign mem_MPORT_211_mask = 1'h1;
  assign mem_MPORT_211_en = reset;
  assign mem_MPORT_212_data = 2'h0;
  assign mem_MPORT_212_addr = 9'hd4;
  assign mem_MPORT_212_mask = 1'h1;
  assign mem_MPORT_212_en = reset;
  assign mem_MPORT_213_data = 2'h0;
  assign mem_MPORT_213_addr = 9'hd5;
  assign mem_MPORT_213_mask = 1'h1;
  assign mem_MPORT_213_en = reset;
  assign mem_MPORT_214_data = 2'h0;
  assign mem_MPORT_214_addr = 9'hd6;
  assign mem_MPORT_214_mask = 1'h1;
  assign mem_MPORT_214_en = reset;
  assign mem_MPORT_215_data = 2'h0;
  assign mem_MPORT_215_addr = 9'hd7;
  assign mem_MPORT_215_mask = 1'h1;
  assign mem_MPORT_215_en = reset;
  assign mem_MPORT_216_data = 2'h0;
  assign mem_MPORT_216_addr = 9'hd8;
  assign mem_MPORT_216_mask = 1'h1;
  assign mem_MPORT_216_en = reset;
  assign mem_MPORT_217_data = 2'h0;
  assign mem_MPORT_217_addr = 9'hd9;
  assign mem_MPORT_217_mask = 1'h1;
  assign mem_MPORT_217_en = reset;
  assign mem_MPORT_218_data = 2'h0;
  assign mem_MPORT_218_addr = 9'hda;
  assign mem_MPORT_218_mask = 1'h1;
  assign mem_MPORT_218_en = reset;
  assign mem_MPORT_219_data = 2'h0;
  assign mem_MPORT_219_addr = 9'hdb;
  assign mem_MPORT_219_mask = 1'h1;
  assign mem_MPORT_219_en = reset;
  assign mem_MPORT_220_data = 2'h0;
  assign mem_MPORT_220_addr = 9'hdc;
  assign mem_MPORT_220_mask = 1'h1;
  assign mem_MPORT_220_en = reset;
  assign mem_MPORT_221_data = 2'h0;
  assign mem_MPORT_221_addr = 9'hdd;
  assign mem_MPORT_221_mask = 1'h1;
  assign mem_MPORT_221_en = reset;
  assign mem_MPORT_222_data = 2'h0;
  assign mem_MPORT_222_addr = 9'hde;
  assign mem_MPORT_222_mask = 1'h1;
  assign mem_MPORT_222_en = reset;
  assign mem_MPORT_223_data = 2'h0;
  assign mem_MPORT_223_addr = 9'hdf;
  assign mem_MPORT_223_mask = 1'h1;
  assign mem_MPORT_223_en = reset;
  assign mem_MPORT_224_data = 2'h0;
  assign mem_MPORT_224_addr = 9'he0;
  assign mem_MPORT_224_mask = 1'h1;
  assign mem_MPORT_224_en = reset;
  assign mem_MPORT_225_data = 2'h0;
  assign mem_MPORT_225_addr = 9'he1;
  assign mem_MPORT_225_mask = 1'h1;
  assign mem_MPORT_225_en = reset;
  assign mem_MPORT_226_data = 2'h0;
  assign mem_MPORT_226_addr = 9'he2;
  assign mem_MPORT_226_mask = 1'h1;
  assign mem_MPORT_226_en = reset;
  assign mem_MPORT_227_data = 2'h0;
  assign mem_MPORT_227_addr = 9'he3;
  assign mem_MPORT_227_mask = 1'h1;
  assign mem_MPORT_227_en = reset;
  assign mem_MPORT_228_data = 2'h0;
  assign mem_MPORT_228_addr = 9'he4;
  assign mem_MPORT_228_mask = 1'h1;
  assign mem_MPORT_228_en = reset;
  assign mem_MPORT_229_data = 2'h0;
  assign mem_MPORT_229_addr = 9'he5;
  assign mem_MPORT_229_mask = 1'h1;
  assign mem_MPORT_229_en = reset;
  assign mem_MPORT_230_data = 2'h0;
  assign mem_MPORT_230_addr = 9'he6;
  assign mem_MPORT_230_mask = 1'h1;
  assign mem_MPORT_230_en = reset;
  assign mem_MPORT_231_data = 2'h0;
  assign mem_MPORT_231_addr = 9'he7;
  assign mem_MPORT_231_mask = 1'h1;
  assign mem_MPORT_231_en = reset;
  assign mem_MPORT_232_data = 2'h0;
  assign mem_MPORT_232_addr = 9'he8;
  assign mem_MPORT_232_mask = 1'h1;
  assign mem_MPORT_232_en = reset;
  assign mem_MPORT_233_data = 2'h0;
  assign mem_MPORT_233_addr = 9'he9;
  assign mem_MPORT_233_mask = 1'h1;
  assign mem_MPORT_233_en = reset;
  assign mem_MPORT_234_data = 2'h0;
  assign mem_MPORT_234_addr = 9'hea;
  assign mem_MPORT_234_mask = 1'h1;
  assign mem_MPORT_234_en = reset;
  assign mem_MPORT_235_data = 2'h0;
  assign mem_MPORT_235_addr = 9'heb;
  assign mem_MPORT_235_mask = 1'h1;
  assign mem_MPORT_235_en = reset;
  assign mem_MPORT_236_data = 2'h0;
  assign mem_MPORT_236_addr = 9'hec;
  assign mem_MPORT_236_mask = 1'h1;
  assign mem_MPORT_236_en = reset;
  assign mem_MPORT_237_data = 2'h0;
  assign mem_MPORT_237_addr = 9'hed;
  assign mem_MPORT_237_mask = 1'h1;
  assign mem_MPORT_237_en = reset;
  assign mem_MPORT_238_data = 2'h0;
  assign mem_MPORT_238_addr = 9'hee;
  assign mem_MPORT_238_mask = 1'h1;
  assign mem_MPORT_238_en = reset;
  assign mem_MPORT_239_data = 2'h0;
  assign mem_MPORT_239_addr = 9'hef;
  assign mem_MPORT_239_mask = 1'h1;
  assign mem_MPORT_239_en = reset;
  assign mem_MPORT_240_data = 2'h0;
  assign mem_MPORT_240_addr = 9'hf0;
  assign mem_MPORT_240_mask = 1'h1;
  assign mem_MPORT_240_en = reset;
  assign mem_MPORT_241_data = 2'h0;
  assign mem_MPORT_241_addr = 9'hf1;
  assign mem_MPORT_241_mask = 1'h1;
  assign mem_MPORT_241_en = reset;
  assign mem_MPORT_242_data = 2'h0;
  assign mem_MPORT_242_addr = 9'hf2;
  assign mem_MPORT_242_mask = 1'h1;
  assign mem_MPORT_242_en = reset;
  assign mem_MPORT_243_data = 2'h0;
  assign mem_MPORT_243_addr = 9'hf3;
  assign mem_MPORT_243_mask = 1'h1;
  assign mem_MPORT_243_en = reset;
  assign mem_MPORT_244_data = 2'h0;
  assign mem_MPORT_244_addr = 9'hf4;
  assign mem_MPORT_244_mask = 1'h1;
  assign mem_MPORT_244_en = reset;
  assign mem_MPORT_245_data = 2'h0;
  assign mem_MPORT_245_addr = 9'hf5;
  assign mem_MPORT_245_mask = 1'h1;
  assign mem_MPORT_245_en = reset;
  assign mem_MPORT_246_data = 2'h0;
  assign mem_MPORT_246_addr = 9'hf6;
  assign mem_MPORT_246_mask = 1'h1;
  assign mem_MPORT_246_en = reset;
  assign mem_MPORT_247_data = 2'h0;
  assign mem_MPORT_247_addr = 9'hf7;
  assign mem_MPORT_247_mask = 1'h1;
  assign mem_MPORT_247_en = reset;
  assign mem_MPORT_248_data = 2'h0;
  assign mem_MPORT_248_addr = 9'hf8;
  assign mem_MPORT_248_mask = 1'h1;
  assign mem_MPORT_248_en = reset;
  assign mem_MPORT_249_data = 2'h0;
  assign mem_MPORT_249_addr = 9'hf9;
  assign mem_MPORT_249_mask = 1'h1;
  assign mem_MPORT_249_en = reset;
  assign mem_MPORT_250_data = 2'h0;
  assign mem_MPORT_250_addr = 9'hfa;
  assign mem_MPORT_250_mask = 1'h1;
  assign mem_MPORT_250_en = reset;
  assign mem_MPORT_251_data = 2'h0;
  assign mem_MPORT_251_addr = 9'hfb;
  assign mem_MPORT_251_mask = 1'h1;
  assign mem_MPORT_251_en = reset;
  assign mem_MPORT_252_data = 2'h0;
  assign mem_MPORT_252_addr = 9'hfc;
  assign mem_MPORT_252_mask = 1'h1;
  assign mem_MPORT_252_en = reset;
  assign mem_MPORT_253_data = 2'h0;
  assign mem_MPORT_253_addr = 9'hfd;
  assign mem_MPORT_253_mask = 1'h1;
  assign mem_MPORT_253_en = reset;
  assign mem_MPORT_254_data = 2'h0;
  assign mem_MPORT_254_addr = 9'hfe;
  assign mem_MPORT_254_mask = 1'h1;
  assign mem_MPORT_254_en = reset;
  assign mem_MPORT_255_data = 2'h0;
  assign mem_MPORT_255_addr = 9'hff;
  assign mem_MPORT_255_mask = 1'h1;
  assign mem_MPORT_255_en = reset;
  assign mem_MPORT_256_data = 2'h0;
  assign mem_MPORT_256_addr = 9'h100;
  assign mem_MPORT_256_mask = 1'h1;
  assign mem_MPORT_256_en = reset;
  assign mem_MPORT_257_data = 2'h0;
  assign mem_MPORT_257_addr = 9'h101;
  assign mem_MPORT_257_mask = 1'h1;
  assign mem_MPORT_257_en = reset;
  assign mem_MPORT_258_data = 2'h0;
  assign mem_MPORT_258_addr = 9'h102;
  assign mem_MPORT_258_mask = 1'h1;
  assign mem_MPORT_258_en = reset;
  assign mem_MPORT_259_data = 2'h0;
  assign mem_MPORT_259_addr = 9'h103;
  assign mem_MPORT_259_mask = 1'h1;
  assign mem_MPORT_259_en = reset;
  assign mem_MPORT_260_data = 2'h0;
  assign mem_MPORT_260_addr = 9'h104;
  assign mem_MPORT_260_mask = 1'h1;
  assign mem_MPORT_260_en = reset;
  assign mem_MPORT_261_data = 2'h0;
  assign mem_MPORT_261_addr = 9'h105;
  assign mem_MPORT_261_mask = 1'h1;
  assign mem_MPORT_261_en = reset;
  assign mem_MPORT_262_data = 2'h0;
  assign mem_MPORT_262_addr = 9'h106;
  assign mem_MPORT_262_mask = 1'h1;
  assign mem_MPORT_262_en = reset;
  assign mem_MPORT_263_data = 2'h0;
  assign mem_MPORT_263_addr = 9'h107;
  assign mem_MPORT_263_mask = 1'h1;
  assign mem_MPORT_263_en = reset;
  assign mem_MPORT_264_data = 2'h0;
  assign mem_MPORT_264_addr = 9'h108;
  assign mem_MPORT_264_mask = 1'h1;
  assign mem_MPORT_264_en = reset;
  assign mem_MPORT_265_data = 2'h0;
  assign mem_MPORT_265_addr = 9'h109;
  assign mem_MPORT_265_mask = 1'h1;
  assign mem_MPORT_265_en = reset;
  assign mem_MPORT_266_data = 2'h0;
  assign mem_MPORT_266_addr = 9'h10a;
  assign mem_MPORT_266_mask = 1'h1;
  assign mem_MPORT_266_en = reset;
  assign mem_MPORT_267_data = 2'h0;
  assign mem_MPORT_267_addr = 9'h10b;
  assign mem_MPORT_267_mask = 1'h1;
  assign mem_MPORT_267_en = reset;
  assign mem_MPORT_268_data = 2'h0;
  assign mem_MPORT_268_addr = 9'h10c;
  assign mem_MPORT_268_mask = 1'h1;
  assign mem_MPORT_268_en = reset;
  assign mem_MPORT_269_data = 2'h0;
  assign mem_MPORT_269_addr = 9'h10d;
  assign mem_MPORT_269_mask = 1'h1;
  assign mem_MPORT_269_en = reset;
  assign mem_MPORT_270_data = 2'h0;
  assign mem_MPORT_270_addr = 9'h10e;
  assign mem_MPORT_270_mask = 1'h1;
  assign mem_MPORT_270_en = reset;
  assign mem_MPORT_271_data = 2'h0;
  assign mem_MPORT_271_addr = 9'h10f;
  assign mem_MPORT_271_mask = 1'h1;
  assign mem_MPORT_271_en = reset;
  assign mem_MPORT_272_data = 2'h0;
  assign mem_MPORT_272_addr = 9'h110;
  assign mem_MPORT_272_mask = 1'h1;
  assign mem_MPORT_272_en = reset;
  assign mem_MPORT_273_data = 2'h0;
  assign mem_MPORT_273_addr = 9'h111;
  assign mem_MPORT_273_mask = 1'h1;
  assign mem_MPORT_273_en = reset;
  assign mem_MPORT_274_data = 2'h0;
  assign mem_MPORT_274_addr = 9'h112;
  assign mem_MPORT_274_mask = 1'h1;
  assign mem_MPORT_274_en = reset;
  assign mem_MPORT_275_data = 2'h0;
  assign mem_MPORT_275_addr = 9'h113;
  assign mem_MPORT_275_mask = 1'h1;
  assign mem_MPORT_275_en = reset;
  assign mem_MPORT_276_data = 2'h0;
  assign mem_MPORT_276_addr = 9'h114;
  assign mem_MPORT_276_mask = 1'h1;
  assign mem_MPORT_276_en = reset;
  assign mem_MPORT_277_data = 2'h0;
  assign mem_MPORT_277_addr = 9'h115;
  assign mem_MPORT_277_mask = 1'h1;
  assign mem_MPORT_277_en = reset;
  assign mem_MPORT_278_data = 2'h0;
  assign mem_MPORT_278_addr = 9'h116;
  assign mem_MPORT_278_mask = 1'h1;
  assign mem_MPORT_278_en = reset;
  assign mem_MPORT_279_data = 2'h0;
  assign mem_MPORT_279_addr = 9'h117;
  assign mem_MPORT_279_mask = 1'h1;
  assign mem_MPORT_279_en = reset;
  assign mem_MPORT_280_data = 2'h0;
  assign mem_MPORT_280_addr = 9'h118;
  assign mem_MPORT_280_mask = 1'h1;
  assign mem_MPORT_280_en = reset;
  assign mem_MPORT_281_data = 2'h0;
  assign mem_MPORT_281_addr = 9'h119;
  assign mem_MPORT_281_mask = 1'h1;
  assign mem_MPORT_281_en = reset;
  assign mem_MPORT_282_data = 2'h0;
  assign mem_MPORT_282_addr = 9'h11a;
  assign mem_MPORT_282_mask = 1'h1;
  assign mem_MPORT_282_en = reset;
  assign mem_MPORT_283_data = 2'h0;
  assign mem_MPORT_283_addr = 9'h11b;
  assign mem_MPORT_283_mask = 1'h1;
  assign mem_MPORT_283_en = reset;
  assign mem_MPORT_284_data = 2'h0;
  assign mem_MPORT_284_addr = 9'h11c;
  assign mem_MPORT_284_mask = 1'h1;
  assign mem_MPORT_284_en = reset;
  assign mem_MPORT_285_data = 2'h0;
  assign mem_MPORT_285_addr = 9'h11d;
  assign mem_MPORT_285_mask = 1'h1;
  assign mem_MPORT_285_en = reset;
  assign mem_MPORT_286_data = 2'h0;
  assign mem_MPORT_286_addr = 9'h11e;
  assign mem_MPORT_286_mask = 1'h1;
  assign mem_MPORT_286_en = reset;
  assign mem_MPORT_287_data = 2'h0;
  assign mem_MPORT_287_addr = 9'h11f;
  assign mem_MPORT_287_mask = 1'h1;
  assign mem_MPORT_287_en = reset;
  assign mem_MPORT_288_data = 2'h0;
  assign mem_MPORT_288_addr = 9'h120;
  assign mem_MPORT_288_mask = 1'h1;
  assign mem_MPORT_288_en = reset;
  assign mem_MPORT_289_data = 2'h0;
  assign mem_MPORT_289_addr = 9'h121;
  assign mem_MPORT_289_mask = 1'h1;
  assign mem_MPORT_289_en = reset;
  assign mem_MPORT_290_data = 2'h0;
  assign mem_MPORT_290_addr = 9'h122;
  assign mem_MPORT_290_mask = 1'h1;
  assign mem_MPORT_290_en = reset;
  assign mem_MPORT_291_data = 2'h0;
  assign mem_MPORT_291_addr = 9'h123;
  assign mem_MPORT_291_mask = 1'h1;
  assign mem_MPORT_291_en = reset;
  assign mem_MPORT_292_data = 2'h0;
  assign mem_MPORT_292_addr = 9'h124;
  assign mem_MPORT_292_mask = 1'h1;
  assign mem_MPORT_292_en = reset;
  assign mem_MPORT_293_data = 2'h0;
  assign mem_MPORT_293_addr = 9'h125;
  assign mem_MPORT_293_mask = 1'h1;
  assign mem_MPORT_293_en = reset;
  assign mem_MPORT_294_data = 2'h0;
  assign mem_MPORT_294_addr = 9'h126;
  assign mem_MPORT_294_mask = 1'h1;
  assign mem_MPORT_294_en = reset;
  assign mem_MPORT_295_data = 2'h0;
  assign mem_MPORT_295_addr = 9'h127;
  assign mem_MPORT_295_mask = 1'h1;
  assign mem_MPORT_295_en = reset;
  assign mem_MPORT_296_data = 2'h0;
  assign mem_MPORT_296_addr = 9'h128;
  assign mem_MPORT_296_mask = 1'h1;
  assign mem_MPORT_296_en = reset;
  assign mem_MPORT_297_data = 2'h0;
  assign mem_MPORT_297_addr = 9'h129;
  assign mem_MPORT_297_mask = 1'h1;
  assign mem_MPORT_297_en = reset;
  assign mem_MPORT_298_data = 2'h0;
  assign mem_MPORT_298_addr = 9'h12a;
  assign mem_MPORT_298_mask = 1'h1;
  assign mem_MPORT_298_en = reset;
  assign mem_MPORT_299_data = 2'h0;
  assign mem_MPORT_299_addr = 9'h12b;
  assign mem_MPORT_299_mask = 1'h1;
  assign mem_MPORT_299_en = reset;
  assign mem_MPORT_300_data = 2'h0;
  assign mem_MPORT_300_addr = 9'h12c;
  assign mem_MPORT_300_mask = 1'h1;
  assign mem_MPORT_300_en = reset;
  assign mem_MPORT_301_data = 2'h0;
  assign mem_MPORT_301_addr = 9'h12d;
  assign mem_MPORT_301_mask = 1'h1;
  assign mem_MPORT_301_en = reset;
  assign mem_MPORT_302_data = 2'h0;
  assign mem_MPORT_302_addr = 9'h12e;
  assign mem_MPORT_302_mask = 1'h1;
  assign mem_MPORT_302_en = reset;
  assign mem_MPORT_303_data = 2'h0;
  assign mem_MPORT_303_addr = 9'h12f;
  assign mem_MPORT_303_mask = 1'h1;
  assign mem_MPORT_303_en = reset;
  assign mem_MPORT_304_data = 2'h0;
  assign mem_MPORT_304_addr = 9'h130;
  assign mem_MPORT_304_mask = 1'h1;
  assign mem_MPORT_304_en = reset;
  assign mem_MPORT_305_data = 2'h0;
  assign mem_MPORT_305_addr = 9'h131;
  assign mem_MPORT_305_mask = 1'h1;
  assign mem_MPORT_305_en = reset;
  assign mem_MPORT_306_data = 2'h0;
  assign mem_MPORT_306_addr = 9'h132;
  assign mem_MPORT_306_mask = 1'h1;
  assign mem_MPORT_306_en = reset;
  assign mem_MPORT_307_data = 2'h0;
  assign mem_MPORT_307_addr = 9'h133;
  assign mem_MPORT_307_mask = 1'h1;
  assign mem_MPORT_307_en = reset;
  assign mem_MPORT_308_data = 2'h0;
  assign mem_MPORT_308_addr = 9'h134;
  assign mem_MPORT_308_mask = 1'h1;
  assign mem_MPORT_308_en = reset;
  assign mem_MPORT_309_data = 2'h0;
  assign mem_MPORT_309_addr = 9'h135;
  assign mem_MPORT_309_mask = 1'h1;
  assign mem_MPORT_309_en = reset;
  assign mem_MPORT_310_data = 2'h0;
  assign mem_MPORT_310_addr = 9'h136;
  assign mem_MPORT_310_mask = 1'h1;
  assign mem_MPORT_310_en = reset;
  assign mem_MPORT_311_data = 2'h0;
  assign mem_MPORT_311_addr = 9'h137;
  assign mem_MPORT_311_mask = 1'h1;
  assign mem_MPORT_311_en = reset;
  assign mem_MPORT_312_data = 2'h0;
  assign mem_MPORT_312_addr = 9'h138;
  assign mem_MPORT_312_mask = 1'h1;
  assign mem_MPORT_312_en = reset;
  assign mem_MPORT_313_data = 2'h0;
  assign mem_MPORT_313_addr = 9'h139;
  assign mem_MPORT_313_mask = 1'h1;
  assign mem_MPORT_313_en = reset;
  assign mem_MPORT_314_data = 2'h0;
  assign mem_MPORT_314_addr = 9'h13a;
  assign mem_MPORT_314_mask = 1'h1;
  assign mem_MPORT_314_en = reset;
  assign mem_MPORT_315_data = 2'h0;
  assign mem_MPORT_315_addr = 9'h13b;
  assign mem_MPORT_315_mask = 1'h1;
  assign mem_MPORT_315_en = reset;
  assign mem_MPORT_316_data = 2'h0;
  assign mem_MPORT_316_addr = 9'h13c;
  assign mem_MPORT_316_mask = 1'h1;
  assign mem_MPORT_316_en = reset;
  assign mem_MPORT_317_data = 2'h0;
  assign mem_MPORT_317_addr = 9'h13d;
  assign mem_MPORT_317_mask = 1'h1;
  assign mem_MPORT_317_en = reset;
  assign mem_MPORT_318_data = 2'h0;
  assign mem_MPORT_318_addr = 9'h13e;
  assign mem_MPORT_318_mask = 1'h1;
  assign mem_MPORT_318_en = reset;
  assign mem_MPORT_319_data = 2'h0;
  assign mem_MPORT_319_addr = 9'h13f;
  assign mem_MPORT_319_mask = 1'h1;
  assign mem_MPORT_319_en = reset;
  assign mem_MPORT_320_data = 2'h0;
  assign mem_MPORT_320_addr = 9'h140;
  assign mem_MPORT_320_mask = 1'h1;
  assign mem_MPORT_320_en = reset;
  assign mem_MPORT_321_data = 2'h0;
  assign mem_MPORT_321_addr = 9'h141;
  assign mem_MPORT_321_mask = 1'h1;
  assign mem_MPORT_321_en = reset;
  assign mem_MPORT_322_data = 2'h0;
  assign mem_MPORT_322_addr = 9'h142;
  assign mem_MPORT_322_mask = 1'h1;
  assign mem_MPORT_322_en = reset;
  assign mem_MPORT_323_data = 2'h0;
  assign mem_MPORT_323_addr = 9'h143;
  assign mem_MPORT_323_mask = 1'h1;
  assign mem_MPORT_323_en = reset;
  assign mem_MPORT_324_data = 2'h0;
  assign mem_MPORT_324_addr = 9'h144;
  assign mem_MPORT_324_mask = 1'h1;
  assign mem_MPORT_324_en = reset;
  assign mem_MPORT_325_data = 2'h0;
  assign mem_MPORT_325_addr = 9'h145;
  assign mem_MPORT_325_mask = 1'h1;
  assign mem_MPORT_325_en = reset;
  assign mem_MPORT_326_data = 2'h0;
  assign mem_MPORT_326_addr = 9'h146;
  assign mem_MPORT_326_mask = 1'h1;
  assign mem_MPORT_326_en = reset;
  assign mem_MPORT_327_data = 2'h0;
  assign mem_MPORT_327_addr = 9'h147;
  assign mem_MPORT_327_mask = 1'h1;
  assign mem_MPORT_327_en = reset;
  assign mem_MPORT_328_data = 2'h0;
  assign mem_MPORT_328_addr = 9'h148;
  assign mem_MPORT_328_mask = 1'h1;
  assign mem_MPORT_328_en = reset;
  assign mem_MPORT_329_data = 2'h0;
  assign mem_MPORT_329_addr = 9'h149;
  assign mem_MPORT_329_mask = 1'h1;
  assign mem_MPORT_329_en = reset;
  assign mem_MPORT_330_data = 2'h0;
  assign mem_MPORT_330_addr = 9'h14a;
  assign mem_MPORT_330_mask = 1'h1;
  assign mem_MPORT_330_en = reset;
  assign mem_MPORT_331_data = 2'h0;
  assign mem_MPORT_331_addr = 9'h14b;
  assign mem_MPORT_331_mask = 1'h1;
  assign mem_MPORT_331_en = reset;
  assign mem_MPORT_332_data = 2'h0;
  assign mem_MPORT_332_addr = 9'h14c;
  assign mem_MPORT_332_mask = 1'h1;
  assign mem_MPORT_332_en = reset;
  assign mem_MPORT_333_data = 2'h0;
  assign mem_MPORT_333_addr = 9'h14d;
  assign mem_MPORT_333_mask = 1'h1;
  assign mem_MPORT_333_en = reset;
  assign mem_MPORT_334_data = 2'h0;
  assign mem_MPORT_334_addr = 9'h14e;
  assign mem_MPORT_334_mask = 1'h1;
  assign mem_MPORT_334_en = reset;
  assign mem_MPORT_335_data = 2'h0;
  assign mem_MPORT_335_addr = 9'h14f;
  assign mem_MPORT_335_mask = 1'h1;
  assign mem_MPORT_335_en = reset;
  assign mem_MPORT_336_data = 2'h0;
  assign mem_MPORT_336_addr = 9'h150;
  assign mem_MPORT_336_mask = 1'h1;
  assign mem_MPORT_336_en = reset;
  assign mem_MPORT_337_data = 2'h0;
  assign mem_MPORT_337_addr = 9'h151;
  assign mem_MPORT_337_mask = 1'h1;
  assign mem_MPORT_337_en = reset;
  assign mem_MPORT_338_data = 2'h0;
  assign mem_MPORT_338_addr = 9'h152;
  assign mem_MPORT_338_mask = 1'h1;
  assign mem_MPORT_338_en = reset;
  assign mem_MPORT_339_data = 2'h0;
  assign mem_MPORT_339_addr = 9'h153;
  assign mem_MPORT_339_mask = 1'h1;
  assign mem_MPORT_339_en = reset;
  assign mem_MPORT_340_data = 2'h0;
  assign mem_MPORT_340_addr = 9'h154;
  assign mem_MPORT_340_mask = 1'h1;
  assign mem_MPORT_340_en = reset;
  assign mem_MPORT_341_data = 2'h0;
  assign mem_MPORT_341_addr = 9'h155;
  assign mem_MPORT_341_mask = 1'h1;
  assign mem_MPORT_341_en = reset;
  assign mem_MPORT_342_data = 2'h0;
  assign mem_MPORT_342_addr = 9'h156;
  assign mem_MPORT_342_mask = 1'h1;
  assign mem_MPORT_342_en = reset;
  assign mem_MPORT_343_data = 2'h0;
  assign mem_MPORT_343_addr = 9'h157;
  assign mem_MPORT_343_mask = 1'h1;
  assign mem_MPORT_343_en = reset;
  assign mem_MPORT_344_data = 2'h0;
  assign mem_MPORT_344_addr = 9'h158;
  assign mem_MPORT_344_mask = 1'h1;
  assign mem_MPORT_344_en = reset;
  assign mem_MPORT_345_data = 2'h0;
  assign mem_MPORT_345_addr = 9'h159;
  assign mem_MPORT_345_mask = 1'h1;
  assign mem_MPORT_345_en = reset;
  assign mem_MPORT_346_data = 2'h0;
  assign mem_MPORT_346_addr = 9'h15a;
  assign mem_MPORT_346_mask = 1'h1;
  assign mem_MPORT_346_en = reset;
  assign mem_MPORT_347_data = 2'h0;
  assign mem_MPORT_347_addr = 9'h15b;
  assign mem_MPORT_347_mask = 1'h1;
  assign mem_MPORT_347_en = reset;
  assign mem_MPORT_348_data = 2'h0;
  assign mem_MPORT_348_addr = 9'h15c;
  assign mem_MPORT_348_mask = 1'h1;
  assign mem_MPORT_348_en = reset;
  assign mem_MPORT_349_data = 2'h0;
  assign mem_MPORT_349_addr = 9'h15d;
  assign mem_MPORT_349_mask = 1'h1;
  assign mem_MPORT_349_en = reset;
  assign mem_MPORT_350_data = 2'h0;
  assign mem_MPORT_350_addr = 9'h15e;
  assign mem_MPORT_350_mask = 1'h1;
  assign mem_MPORT_350_en = reset;
  assign mem_MPORT_351_data = 2'h0;
  assign mem_MPORT_351_addr = 9'h15f;
  assign mem_MPORT_351_mask = 1'h1;
  assign mem_MPORT_351_en = reset;
  assign mem_MPORT_352_data = 2'h0;
  assign mem_MPORT_352_addr = 9'h160;
  assign mem_MPORT_352_mask = 1'h1;
  assign mem_MPORT_352_en = reset;
  assign mem_MPORT_353_data = 2'h0;
  assign mem_MPORT_353_addr = 9'h161;
  assign mem_MPORT_353_mask = 1'h1;
  assign mem_MPORT_353_en = reset;
  assign mem_MPORT_354_data = 2'h0;
  assign mem_MPORT_354_addr = 9'h162;
  assign mem_MPORT_354_mask = 1'h1;
  assign mem_MPORT_354_en = reset;
  assign mem_MPORT_355_data = 2'h0;
  assign mem_MPORT_355_addr = 9'h163;
  assign mem_MPORT_355_mask = 1'h1;
  assign mem_MPORT_355_en = reset;
  assign mem_MPORT_356_data = 2'h0;
  assign mem_MPORT_356_addr = 9'h164;
  assign mem_MPORT_356_mask = 1'h1;
  assign mem_MPORT_356_en = reset;
  assign mem_MPORT_357_data = 2'h0;
  assign mem_MPORT_357_addr = 9'h165;
  assign mem_MPORT_357_mask = 1'h1;
  assign mem_MPORT_357_en = reset;
  assign mem_MPORT_358_data = 2'h0;
  assign mem_MPORT_358_addr = 9'h166;
  assign mem_MPORT_358_mask = 1'h1;
  assign mem_MPORT_358_en = reset;
  assign mem_MPORT_359_data = 2'h0;
  assign mem_MPORT_359_addr = 9'h167;
  assign mem_MPORT_359_mask = 1'h1;
  assign mem_MPORT_359_en = reset;
  assign mem_MPORT_360_data = 2'h0;
  assign mem_MPORT_360_addr = 9'h168;
  assign mem_MPORT_360_mask = 1'h1;
  assign mem_MPORT_360_en = reset;
  assign mem_MPORT_361_data = 2'h0;
  assign mem_MPORT_361_addr = 9'h169;
  assign mem_MPORT_361_mask = 1'h1;
  assign mem_MPORT_361_en = reset;
  assign mem_MPORT_362_data = 2'h0;
  assign mem_MPORT_362_addr = 9'h16a;
  assign mem_MPORT_362_mask = 1'h1;
  assign mem_MPORT_362_en = reset;
  assign mem_MPORT_363_data = 2'h0;
  assign mem_MPORT_363_addr = 9'h16b;
  assign mem_MPORT_363_mask = 1'h1;
  assign mem_MPORT_363_en = reset;
  assign mem_MPORT_364_data = 2'h0;
  assign mem_MPORT_364_addr = 9'h16c;
  assign mem_MPORT_364_mask = 1'h1;
  assign mem_MPORT_364_en = reset;
  assign mem_MPORT_365_data = 2'h0;
  assign mem_MPORT_365_addr = 9'h16d;
  assign mem_MPORT_365_mask = 1'h1;
  assign mem_MPORT_365_en = reset;
  assign mem_MPORT_366_data = 2'h0;
  assign mem_MPORT_366_addr = 9'h16e;
  assign mem_MPORT_366_mask = 1'h1;
  assign mem_MPORT_366_en = reset;
  assign mem_MPORT_367_data = 2'h0;
  assign mem_MPORT_367_addr = 9'h16f;
  assign mem_MPORT_367_mask = 1'h1;
  assign mem_MPORT_367_en = reset;
  assign mem_MPORT_368_data = 2'h0;
  assign mem_MPORT_368_addr = 9'h170;
  assign mem_MPORT_368_mask = 1'h1;
  assign mem_MPORT_368_en = reset;
  assign mem_MPORT_369_data = 2'h0;
  assign mem_MPORT_369_addr = 9'h171;
  assign mem_MPORT_369_mask = 1'h1;
  assign mem_MPORT_369_en = reset;
  assign mem_MPORT_370_data = 2'h0;
  assign mem_MPORT_370_addr = 9'h172;
  assign mem_MPORT_370_mask = 1'h1;
  assign mem_MPORT_370_en = reset;
  assign mem_MPORT_371_data = 2'h0;
  assign mem_MPORT_371_addr = 9'h173;
  assign mem_MPORT_371_mask = 1'h1;
  assign mem_MPORT_371_en = reset;
  assign mem_MPORT_372_data = 2'h0;
  assign mem_MPORT_372_addr = 9'h174;
  assign mem_MPORT_372_mask = 1'h1;
  assign mem_MPORT_372_en = reset;
  assign mem_MPORT_373_data = 2'h0;
  assign mem_MPORT_373_addr = 9'h175;
  assign mem_MPORT_373_mask = 1'h1;
  assign mem_MPORT_373_en = reset;
  assign mem_MPORT_374_data = 2'h0;
  assign mem_MPORT_374_addr = 9'h176;
  assign mem_MPORT_374_mask = 1'h1;
  assign mem_MPORT_374_en = reset;
  assign mem_MPORT_375_data = 2'h0;
  assign mem_MPORT_375_addr = 9'h177;
  assign mem_MPORT_375_mask = 1'h1;
  assign mem_MPORT_375_en = reset;
  assign mem_MPORT_376_data = 2'h0;
  assign mem_MPORT_376_addr = 9'h178;
  assign mem_MPORT_376_mask = 1'h1;
  assign mem_MPORT_376_en = reset;
  assign mem_MPORT_377_data = 2'h0;
  assign mem_MPORT_377_addr = 9'h179;
  assign mem_MPORT_377_mask = 1'h1;
  assign mem_MPORT_377_en = reset;
  assign mem_MPORT_378_data = 2'h0;
  assign mem_MPORT_378_addr = 9'h17a;
  assign mem_MPORT_378_mask = 1'h1;
  assign mem_MPORT_378_en = reset;
  assign mem_MPORT_379_data = 2'h0;
  assign mem_MPORT_379_addr = 9'h17b;
  assign mem_MPORT_379_mask = 1'h1;
  assign mem_MPORT_379_en = reset;
  assign mem_MPORT_380_data = 2'h0;
  assign mem_MPORT_380_addr = 9'h17c;
  assign mem_MPORT_380_mask = 1'h1;
  assign mem_MPORT_380_en = reset;
  assign mem_MPORT_381_data = 2'h0;
  assign mem_MPORT_381_addr = 9'h17d;
  assign mem_MPORT_381_mask = 1'h1;
  assign mem_MPORT_381_en = reset;
  assign mem_MPORT_382_data = 2'h0;
  assign mem_MPORT_382_addr = 9'h17e;
  assign mem_MPORT_382_mask = 1'h1;
  assign mem_MPORT_382_en = reset;
  assign mem_MPORT_383_data = 2'h0;
  assign mem_MPORT_383_addr = 9'h17f;
  assign mem_MPORT_383_mask = 1'h1;
  assign mem_MPORT_383_en = reset;
  assign mem_MPORT_384_data = 2'h0;
  assign mem_MPORT_384_addr = 9'h180;
  assign mem_MPORT_384_mask = 1'h1;
  assign mem_MPORT_384_en = reset;
  assign mem_MPORT_385_data = 2'h0;
  assign mem_MPORT_385_addr = 9'h181;
  assign mem_MPORT_385_mask = 1'h1;
  assign mem_MPORT_385_en = reset;
  assign mem_MPORT_386_data = 2'h0;
  assign mem_MPORT_386_addr = 9'h182;
  assign mem_MPORT_386_mask = 1'h1;
  assign mem_MPORT_386_en = reset;
  assign mem_MPORT_387_data = 2'h0;
  assign mem_MPORT_387_addr = 9'h183;
  assign mem_MPORT_387_mask = 1'h1;
  assign mem_MPORT_387_en = reset;
  assign mem_MPORT_388_data = 2'h0;
  assign mem_MPORT_388_addr = 9'h184;
  assign mem_MPORT_388_mask = 1'h1;
  assign mem_MPORT_388_en = reset;
  assign mem_MPORT_389_data = 2'h0;
  assign mem_MPORT_389_addr = 9'h185;
  assign mem_MPORT_389_mask = 1'h1;
  assign mem_MPORT_389_en = reset;
  assign mem_MPORT_390_data = 2'h0;
  assign mem_MPORT_390_addr = 9'h186;
  assign mem_MPORT_390_mask = 1'h1;
  assign mem_MPORT_390_en = reset;
  assign mem_MPORT_391_data = 2'h0;
  assign mem_MPORT_391_addr = 9'h187;
  assign mem_MPORT_391_mask = 1'h1;
  assign mem_MPORT_391_en = reset;
  assign mem_MPORT_392_data = 2'h0;
  assign mem_MPORT_392_addr = 9'h188;
  assign mem_MPORT_392_mask = 1'h1;
  assign mem_MPORT_392_en = reset;
  assign mem_MPORT_393_data = 2'h0;
  assign mem_MPORT_393_addr = 9'h189;
  assign mem_MPORT_393_mask = 1'h1;
  assign mem_MPORT_393_en = reset;
  assign mem_MPORT_394_data = 2'h0;
  assign mem_MPORT_394_addr = 9'h18a;
  assign mem_MPORT_394_mask = 1'h1;
  assign mem_MPORT_394_en = reset;
  assign mem_MPORT_395_data = 2'h0;
  assign mem_MPORT_395_addr = 9'h18b;
  assign mem_MPORT_395_mask = 1'h1;
  assign mem_MPORT_395_en = reset;
  assign mem_MPORT_396_data = 2'h0;
  assign mem_MPORT_396_addr = 9'h18c;
  assign mem_MPORT_396_mask = 1'h1;
  assign mem_MPORT_396_en = reset;
  assign mem_MPORT_397_data = 2'h0;
  assign mem_MPORT_397_addr = 9'h18d;
  assign mem_MPORT_397_mask = 1'h1;
  assign mem_MPORT_397_en = reset;
  assign mem_MPORT_398_data = 2'h0;
  assign mem_MPORT_398_addr = 9'h18e;
  assign mem_MPORT_398_mask = 1'h1;
  assign mem_MPORT_398_en = reset;
  assign mem_MPORT_399_data = 2'h0;
  assign mem_MPORT_399_addr = 9'h18f;
  assign mem_MPORT_399_mask = 1'h1;
  assign mem_MPORT_399_en = reset;
  assign mem_MPORT_400_data = 2'h0;
  assign mem_MPORT_400_addr = 9'h190;
  assign mem_MPORT_400_mask = 1'h1;
  assign mem_MPORT_400_en = reset;
  assign mem_MPORT_401_data = 2'h0;
  assign mem_MPORT_401_addr = 9'h191;
  assign mem_MPORT_401_mask = 1'h1;
  assign mem_MPORT_401_en = reset;
  assign mem_MPORT_402_data = 2'h0;
  assign mem_MPORT_402_addr = 9'h192;
  assign mem_MPORT_402_mask = 1'h1;
  assign mem_MPORT_402_en = reset;
  assign mem_MPORT_403_data = 2'h0;
  assign mem_MPORT_403_addr = 9'h193;
  assign mem_MPORT_403_mask = 1'h1;
  assign mem_MPORT_403_en = reset;
  assign mem_MPORT_404_data = 2'h0;
  assign mem_MPORT_404_addr = 9'h194;
  assign mem_MPORT_404_mask = 1'h1;
  assign mem_MPORT_404_en = reset;
  assign mem_MPORT_405_data = 2'h0;
  assign mem_MPORT_405_addr = 9'h195;
  assign mem_MPORT_405_mask = 1'h1;
  assign mem_MPORT_405_en = reset;
  assign mem_MPORT_406_data = 2'h0;
  assign mem_MPORT_406_addr = 9'h196;
  assign mem_MPORT_406_mask = 1'h1;
  assign mem_MPORT_406_en = reset;
  assign mem_MPORT_407_data = 2'h0;
  assign mem_MPORT_407_addr = 9'h197;
  assign mem_MPORT_407_mask = 1'h1;
  assign mem_MPORT_407_en = reset;
  assign mem_MPORT_408_data = 2'h0;
  assign mem_MPORT_408_addr = 9'h198;
  assign mem_MPORT_408_mask = 1'h1;
  assign mem_MPORT_408_en = reset;
  assign mem_MPORT_409_data = 2'h0;
  assign mem_MPORT_409_addr = 9'h199;
  assign mem_MPORT_409_mask = 1'h1;
  assign mem_MPORT_409_en = reset;
  assign mem_MPORT_410_data = 2'h0;
  assign mem_MPORT_410_addr = 9'h19a;
  assign mem_MPORT_410_mask = 1'h1;
  assign mem_MPORT_410_en = reset;
  assign mem_MPORT_411_data = 2'h0;
  assign mem_MPORT_411_addr = 9'h19b;
  assign mem_MPORT_411_mask = 1'h1;
  assign mem_MPORT_411_en = reset;
  assign mem_MPORT_412_data = 2'h0;
  assign mem_MPORT_412_addr = 9'h19c;
  assign mem_MPORT_412_mask = 1'h1;
  assign mem_MPORT_412_en = reset;
  assign mem_MPORT_413_data = 2'h0;
  assign mem_MPORT_413_addr = 9'h19d;
  assign mem_MPORT_413_mask = 1'h1;
  assign mem_MPORT_413_en = reset;
  assign mem_MPORT_414_data = 2'h0;
  assign mem_MPORT_414_addr = 9'h19e;
  assign mem_MPORT_414_mask = 1'h1;
  assign mem_MPORT_414_en = reset;
  assign mem_MPORT_415_data = 2'h0;
  assign mem_MPORT_415_addr = 9'h19f;
  assign mem_MPORT_415_mask = 1'h1;
  assign mem_MPORT_415_en = reset;
  assign mem_MPORT_416_data = 2'h0;
  assign mem_MPORT_416_addr = 9'h1a0;
  assign mem_MPORT_416_mask = 1'h1;
  assign mem_MPORT_416_en = reset;
  assign mem_MPORT_417_data = 2'h0;
  assign mem_MPORT_417_addr = 9'h1a1;
  assign mem_MPORT_417_mask = 1'h1;
  assign mem_MPORT_417_en = reset;
  assign mem_MPORT_418_data = 2'h0;
  assign mem_MPORT_418_addr = 9'h1a2;
  assign mem_MPORT_418_mask = 1'h1;
  assign mem_MPORT_418_en = reset;
  assign mem_MPORT_419_data = 2'h0;
  assign mem_MPORT_419_addr = 9'h1a3;
  assign mem_MPORT_419_mask = 1'h1;
  assign mem_MPORT_419_en = reset;
  assign mem_MPORT_420_data = 2'h0;
  assign mem_MPORT_420_addr = 9'h1a4;
  assign mem_MPORT_420_mask = 1'h1;
  assign mem_MPORT_420_en = reset;
  assign mem_MPORT_421_data = 2'h0;
  assign mem_MPORT_421_addr = 9'h1a5;
  assign mem_MPORT_421_mask = 1'h1;
  assign mem_MPORT_421_en = reset;
  assign mem_MPORT_422_data = 2'h0;
  assign mem_MPORT_422_addr = 9'h1a6;
  assign mem_MPORT_422_mask = 1'h1;
  assign mem_MPORT_422_en = reset;
  assign mem_MPORT_423_data = 2'h0;
  assign mem_MPORT_423_addr = 9'h1a7;
  assign mem_MPORT_423_mask = 1'h1;
  assign mem_MPORT_423_en = reset;
  assign mem_MPORT_424_data = 2'h0;
  assign mem_MPORT_424_addr = 9'h1a8;
  assign mem_MPORT_424_mask = 1'h1;
  assign mem_MPORT_424_en = reset;
  assign mem_MPORT_425_data = 2'h0;
  assign mem_MPORT_425_addr = 9'h1a9;
  assign mem_MPORT_425_mask = 1'h1;
  assign mem_MPORT_425_en = reset;
  assign mem_MPORT_426_data = 2'h0;
  assign mem_MPORT_426_addr = 9'h1aa;
  assign mem_MPORT_426_mask = 1'h1;
  assign mem_MPORT_426_en = reset;
  assign mem_MPORT_427_data = 2'h0;
  assign mem_MPORT_427_addr = 9'h1ab;
  assign mem_MPORT_427_mask = 1'h1;
  assign mem_MPORT_427_en = reset;
  assign mem_MPORT_428_data = 2'h0;
  assign mem_MPORT_428_addr = 9'h1ac;
  assign mem_MPORT_428_mask = 1'h1;
  assign mem_MPORT_428_en = reset;
  assign mem_MPORT_429_data = 2'h0;
  assign mem_MPORT_429_addr = 9'h1ad;
  assign mem_MPORT_429_mask = 1'h1;
  assign mem_MPORT_429_en = reset;
  assign mem_MPORT_430_data = 2'h0;
  assign mem_MPORT_430_addr = 9'h1ae;
  assign mem_MPORT_430_mask = 1'h1;
  assign mem_MPORT_430_en = reset;
  assign mem_MPORT_431_data = 2'h0;
  assign mem_MPORT_431_addr = 9'h1af;
  assign mem_MPORT_431_mask = 1'h1;
  assign mem_MPORT_431_en = reset;
  assign mem_MPORT_432_data = 2'h0;
  assign mem_MPORT_432_addr = 9'h1b0;
  assign mem_MPORT_432_mask = 1'h1;
  assign mem_MPORT_432_en = reset;
  assign mem_MPORT_433_data = 2'h0;
  assign mem_MPORT_433_addr = 9'h1b1;
  assign mem_MPORT_433_mask = 1'h1;
  assign mem_MPORT_433_en = reset;
  assign mem_MPORT_434_data = 2'h0;
  assign mem_MPORT_434_addr = 9'h1b2;
  assign mem_MPORT_434_mask = 1'h1;
  assign mem_MPORT_434_en = reset;
  assign mem_MPORT_435_data = 2'h0;
  assign mem_MPORT_435_addr = 9'h1b3;
  assign mem_MPORT_435_mask = 1'h1;
  assign mem_MPORT_435_en = reset;
  assign mem_MPORT_436_data = 2'h0;
  assign mem_MPORT_436_addr = 9'h1b4;
  assign mem_MPORT_436_mask = 1'h1;
  assign mem_MPORT_436_en = reset;
  assign mem_MPORT_437_data = 2'h0;
  assign mem_MPORT_437_addr = 9'h1b5;
  assign mem_MPORT_437_mask = 1'h1;
  assign mem_MPORT_437_en = reset;
  assign mem_MPORT_438_data = 2'h0;
  assign mem_MPORT_438_addr = 9'h1b6;
  assign mem_MPORT_438_mask = 1'h1;
  assign mem_MPORT_438_en = reset;
  assign mem_MPORT_439_data = 2'h0;
  assign mem_MPORT_439_addr = 9'h1b7;
  assign mem_MPORT_439_mask = 1'h1;
  assign mem_MPORT_439_en = reset;
  assign mem_MPORT_440_data = 2'h0;
  assign mem_MPORT_440_addr = 9'h1b8;
  assign mem_MPORT_440_mask = 1'h1;
  assign mem_MPORT_440_en = reset;
  assign mem_MPORT_441_data = 2'h0;
  assign mem_MPORT_441_addr = 9'h1b9;
  assign mem_MPORT_441_mask = 1'h1;
  assign mem_MPORT_441_en = reset;
  assign mem_MPORT_442_data = 2'h0;
  assign mem_MPORT_442_addr = 9'h1ba;
  assign mem_MPORT_442_mask = 1'h1;
  assign mem_MPORT_442_en = reset;
  assign mem_MPORT_443_data = 2'h0;
  assign mem_MPORT_443_addr = 9'h1bb;
  assign mem_MPORT_443_mask = 1'h1;
  assign mem_MPORT_443_en = reset;
  assign mem_MPORT_444_data = 2'h0;
  assign mem_MPORT_444_addr = 9'h1bc;
  assign mem_MPORT_444_mask = 1'h1;
  assign mem_MPORT_444_en = reset;
  assign mem_MPORT_445_data = 2'h0;
  assign mem_MPORT_445_addr = 9'h1bd;
  assign mem_MPORT_445_mask = 1'h1;
  assign mem_MPORT_445_en = reset;
  assign mem_MPORT_446_data = 2'h0;
  assign mem_MPORT_446_addr = 9'h1be;
  assign mem_MPORT_446_mask = 1'h1;
  assign mem_MPORT_446_en = reset;
  assign mem_MPORT_447_data = 2'h0;
  assign mem_MPORT_447_addr = 9'h1bf;
  assign mem_MPORT_447_mask = 1'h1;
  assign mem_MPORT_447_en = reset;
  assign mem_MPORT_448_data = 2'h0;
  assign mem_MPORT_448_addr = 9'h1c0;
  assign mem_MPORT_448_mask = 1'h1;
  assign mem_MPORT_448_en = reset;
  assign mem_MPORT_449_data = 2'h0;
  assign mem_MPORT_449_addr = 9'h1c1;
  assign mem_MPORT_449_mask = 1'h1;
  assign mem_MPORT_449_en = reset;
  assign mem_MPORT_450_data = 2'h0;
  assign mem_MPORT_450_addr = 9'h1c2;
  assign mem_MPORT_450_mask = 1'h1;
  assign mem_MPORT_450_en = reset;
  assign mem_MPORT_451_data = 2'h0;
  assign mem_MPORT_451_addr = 9'h1c3;
  assign mem_MPORT_451_mask = 1'h1;
  assign mem_MPORT_451_en = reset;
  assign mem_MPORT_452_data = 2'h0;
  assign mem_MPORT_452_addr = 9'h1c4;
  assign mem_MPORT_452_mask = 1'h1;
  assign mem_MPORT_452_en = reset;
  assign mem_MPORT_453_data = 2'h0;
  assign mem_MPORT_453_addr = 9'h1c5;
  assign mem_MPORT_453_mask = 1'h1;
  assign mem_MPORT_453_en = reset;
  assign mem_MPORT_454_data = 2'h0;
  assign mem_MPORT_454_addr = 9'h1c6;
  assign mem_MPORT_454_mask = 1'h1;
  assign mem_MPORT_454_en = reset;
  assign mem_MPORT_455_data = 2'h0;
  assign mem_MPORT_455_addr = 9'h1c7;
  assign mem_MPORT_455_mask = 1'h1;
  assign mem_MPORT_455_en = reset;
  assign mem_MPORT_456_data = 2'h0;
  assign mem_MPORT_456_addr = 9'h1c8;
  assign mem_MPORT_456_mask = 1'h1;
  assign mem_MPORT_456_en = reset;
  assign mem_MPORT_457_data = 2'h0;
  assign mem_MPORT_457_addr = 9'h1c9;
  assign mem_MPORT_457_mask = 1'h1;
  assign mem_MPORT_457_en = reset;
  assign mem_MPORT_458_data = 2'h0;
  assign mem_MPORT_458_addr = 9'h1ca;
  assign mem_MPORT_458_mask = 1'h1;
  assign mem_MPORT_458_en = reset;
  assign mem_MPORT_459_data = 2'h0;
  assign mem_MPORT_459_addr = 9'h1cb;
  assign mem_MPORT_459_mask = 1'h1;
  assign mem_MPORT_459_en = reset;
  assign mem_MPORT_460_data = 2'h0;
  assign mem_MPORT_460_addr = 9'h1cc;
  assign mem_MPORT_460_mask = 1'h1;
  assign mem_MPORT_460_en = reset;
  assign mem_MPORT_461_data = 2'h0;
  assign mem_MPORT_461_addr = 9'h1cd;
  assign mem_MPORT_461_mask = 1'h1;
  assign mem_MPORT_461_en = reset;
  assign mem_MPORT_462_data = 2'h0;
  assign mem_MPORT_462_addr = 9'h1ce;
  assign mem_MPORT_462_mask = 1'h1;
  assign mem_MPORT_462_en = reset;
  assign mem_MPORT_463_data = 2'h0;
  assign mem_MPORT_463_addr = 9'h1cf;
  assign mem_MPORT_463_mask = 1'h1;
  assign mem_MPORT_463_en = reset;
  assign mem_MPORT_464_data = 2'h0;
  assign mem_MPORT_464_addr = 9'h1d0;
  assign mem_MPORT_464_mask = 1'h1;
  assign mem_MPORT_464_en = reset;
  assign mem_MPORT_465_data = 2'h0;
  assign mem_MPORT_465_addr = 9'h1d1;
  assign mem_MPORT_465_mask = 1'h1;
  assign mem_MPORT_465_en = reset;
  assign mem_MPORT_466_data = 2'h0;
  assign mem_MPORT_466_addr = 9'h1d2;
  assign mem_MPORT_466_mask = 1'h1;
  assign mem_MPORT_466_en = reset;
  assign mem_MPORT_467_data = 2'h0;
  assign mem_MPORT_467_addr = 9'h1d3;
  assign mem_MPORT_467_mask = 1'h1;
  assign mem_MPORT_467_en = reset;
  assign mem_MPORT_468_data = 2'h0;
  assign mem_MPORT_468_addr = 9'h1d4;
  assign mem_MPORT_468_mask = 1'h1;
  assign mem_MPORT_468_en = reset;
  assign mem_MPORT_469_data = 2'h0;
  assign mem_MPORT_469_addr = 9'h1d5;
  assign mem_MPORT_469_mask = 1'h1;
  assign mem_MPORT_469_en = reset;
  assign mem_MPORT_470_data = 2'h0;
  assign mem_MPORT_470_addr = 9'h1d6;
  assign mem_MPORT_470_mask = 1'h1;
  assign mem_MPORT_470_en = reset;
  assign mem_MPORT_471_data = 2'h0;
  assign mem_MPORT_471_addr = 9'h1d7;
  assign mem_MPORT_471_mask = 1'h1;
  assign mem_MPORT_471_en = reset;
  assign mem_MPORT_472_data = 2'h0;
  assign mem_MPORT_472_addr = 9'h1d8;
  assign mem_MPORT_472_mask = 1'h1;
  assign mem_MPORT_472_en = reset;
  assign mem_MPORT_473_data = 2'h0;
  assign mem_MPORT_473_addr = 9'h1d9;
  assign mem_MPORT_473_mask = 1'h1;
  assign mem_MPORT_473_en = reset;
  assign mem_MPORT_474_data = 2'h0;
  assign mem_MPORT_474_addr = 9'h1da;
  assign mem_MPORT_474_mask = 1'h1;
  assign mem_MPORT_474_en = reset;
  assign mem_MPORT_475_data = 2'h0;
  assign mem_MPORT_475_addr = 9'h1db;
  assign mem_MPORT_475_mask = 1'h1;
  assign mem_MPORT_475_en = reset;
  assign mem_MPORT_476_data = 2'h0;
  assign mem_MPORT_476_addr = 9'h1dc;
  assign mem_MPORT_476_mask = 1'h1;
  assign mem_MPORT_476_en = reset;
  assign mem_MPORT_477_data = 2'h0;
  assign mem_MPORT_477_addr = 9'h1dd;
  assign mem_MPORT_477_mask = 1'h1;
  assign mem_MPORT_477_en = reset;
  assign mem_MPORT_478_data = 2'h0;
  assign mem_MPORT_478_addr = 9'h1de;
  assign mem_MPORT_478_mask = 1'h1;
  assign mem_MPORT_478_en = reset;
  assign mem_MPORT_479_data = 2'h0;
  assign mem_MPORT_479_addr = 9'h1df;
  assign mem_MPORT_479_mask = 1'h1;
  assign mem_MPORT_479_en = reset;
  assign mem_MPORT_480_data = 2'h0;
  assign mem_MPORT_480_addr = 9'h1e0;
  assign mem_MPORT_480_mask = 1'h1;
  assign mem_MPORT_480_en = reset;
  assign mem_MPORT_481_data = 2'h0;
  assign mem_MPORT_481_addr = 9'h1e1;
  assign mem_MPORT_481_mask = 1'h1;
  assign mem_MPORT_481_en = reset;
  assign mem_MPORT_482_data = 2'h0;
  assign mem_MPORT_482_addr = 9'h1e2;
  assign mem_MPORT_482_mask = 1'h1;
  assign mem_MPORT_482_en = reset;
  assign mem_MPORT_483_data = 2'h0;
  assign mem_MPORT_483_addr = 9'h1e3;
  assign mem_MPORT_483_mask = 1'h1;
  assign mem_MPORT_483_en = reset;
  assign mem_MPORT_484_data = 2'h0;
  assign mem_MPORT_484_addr = 9'h1e4;
  assign mem_MPORT_484_mask = 1'h1;
  assign mem_MPORT_484_en = reset;
  assign mem_MPORT_485_data = 2'h0;
  assign mem_MPORT_485_addr = 9'h1e5;
  assign mem_MPORT_485_mask = 1'h1;
  assign mem_MPORT_485_en = reset;
  assign mem_MPORT_486_data = 2'h0;
  assign mem_MPORT_486_addr = 9'h1e6;
  assign mem_MPORT_486_mask = 1'h1;
  assign mem_MPORT_486_en = reset;
  assign mem_MPORT_487_data = 2'h0;
  assign mem_MPORT_487_addr = 9'h1e7;
  assign mem_MPORT_487_mask = 1'h1;
  assign mem_MPORT_487_en = reset;
  assign mem_MPORT_488_data = 2'h0;
  assign mem_MPORT_488_addr = 9'h1e8;
  assign mem_MPORT_488_mask = 1'h1;
  assign mem_MPORT_488_en = reset;
  assign mem_MPORT_489_data = 2'h0;
  assign mem_MPORT_489_addr = 9'h1e9;
  assign mem_MPORT_489_mask = 1'h1;
  assign mem_MPORT_489_en = reset;
  assign mem_MPORT_490_data = 2'h0;
  assign mem_MPORT_490_addr = 9'h1ea;
  assign mem_MPORT_490_mask = 1'h1;
  assign mem_MPORT_490_en = reset;
  assign mem_MPORT_491_data = 2'h0;
  assign mem_MPORT_491_addr = 9'h1eb;
  assign mem_MPORT_491_mask = 1'h1;
  assign mem_MPORT_491_en = reset;
  assign mem_MPORT_492_data = 2'h0;
  assign mem_MPORT_492_addr = 9'h1ec;
  assign mem_MPORT_492_mask = 1'h1;
  assign mem_MPORT_492_en = reset;
  assign mem_MPORT_493_data = 2'h0;
  assign mem_MPORT_493_addr = 9'h1ed;
  assign mem_MPORT_493_mask = 1'h1;
  assign mem_MPORT_493_en = reset;
  assign mem_MPORT_494_data = 2'h0;
  assign mem_MPORT_494_addr = 9'h1ee;
  assign mem_MPORT_494_mask = 1'h1;
  assign mem_MPORT_494_en = reset;
  assign mem_MPORT_495_data = 2'h0;
  assign mem_MPORT_495_addr = 9'h1ef;
  assign mem_MPORT_495_mask = 1'h1;
  assign mem_MPORT_495_en = reset;
  assign mem_MPORT_496_data = 2'h0;
  assign mem_MPORT_496_addr = 9'h1f0;
  assign mem_MPORT_496_mask = 1'h1;
  assign mem_MPORT_496_en = reset;
  assign mem_MPORT_497_data = 2'h0;
  assign mem_MPORT_497_addr = 9'h1f1;
  assign mem_MPORT_497_mask = 1'h1;
  assign mem_MPORT_497_en = reset;
  assign mem_MPORT_498_data = 2'h0;
  assign mem_MPORT_498_addr = 9'h1f2;
  assign mem_MPORT_498_mask = 1'h1;
  assign mem_MPORT_498_en = reset;
  assign mem_MPORT_499_data = 2'h0;
  assign mem_MPORT_499_addr = 9'h1f3;
  assign mem_MPORT_499_mask = 1'h1;
  assign mem_MPORT_499_en = reset;
  assign mem_MPORT_500_data = 2'h0;
  assign mem_MPORT_500_addr = 9'h1f4;
  assign mem_MPORT_500_mask = 1'h1;
  assign mem_MPORT_500_en = reset;
  assign mem_MPORT_501_data = 2'h0;
  assign mem_MPORT_501_addr = 9'h1f5;
  assign mem_MPORT_501_mask = 1'h1;
  assign mem_MPORT_501_en = reset;
  assign mem_MPORT_502_data = 2'h0;
  assign mem_MPORT_502_addr = 9'h1f6;
  assign mem_MPORT_502_mask = 1'h1;
  assign mem_MPORT_502_en = reset;
  assign mem_MPORT_503_data = 2'h0;
  assign mem_MPORT_503_addr = 9'h1f7;
  assign mem_MPORT_503_mask = 1'h1;
  assign mem_MPORT_503_en = reset;
  assign mem_MPORT_504_data = 2'h0;
  assign mem_MPORT_504_addr = 9'h1f8;
  assign mem_MPORT_504_mask = 1'h1;
  assign mem_MPORT_504_en = reset;
  assign mem_MPORT_505_data = 2'h0;
  assign mem_MPORT_505_addr = 9'h1f9;
  assign mem_MPORT_505_mask = 1'h1;
  assign mem_MPORT_505_en = reset;
  assign mem_MPORT_506_data = 2'h0;
  assign mem_MPORT_506_addr = 9'h1fa;
  assign mem_MPORT_506_mask = 1'h1;
  assign mem_MPORT_506_en = reset;
  assign mem_MPORT_507_data = 2'h0;
  assign mem_MPORT_507_addr = 9'h1fb;
  assign mem_MPORT_507_mask = 1'h1;
  assign mem_MPORT_507_en = reset;
  assign mem_MPORT_508_data = 2'h0;
  assign mem_MPORT_508_addr = 9'h1fc;
  assign mem_MPORT_508_mask = 1'h1;
  assign mem_MPORT_508_en = reset;
  assign mem_MPORT_509_data = 2'h0;
  assign mem_MPORT_509_addr = 9'h1fd;
  assign mem_MPORT_509_mask = 1'h1;
  assign mem_MPORT_509_en = reset;
  assign mem_MPORT_510_data = 2'h0;
  assign mem_MPORT_510_addr = 9'h1fe;
  assign mem_MPORT_510_mask = 1'h1;
  assign mem_MPORT_510_en = reset;
  assign mem_MPORT_511_data = 2'h0;
  assign mem_MPORT_511_addr = 9'h1ff;
  assign mem_MPORT_511_mask = 1'h1;
  assign mem_MPORT_511_en = reset;
  assign mem_MPORT_512_data = io_w_data;
  assign mem_MPORT_512_addr = io_w_addr;
  assign mem_MPORT_512_mask = 1'h1;
  assign mem_MPORT_512_en = io_w_en;
  assign io_r_data = io_w_en & readConflict ? io_w_data : mem_io_r_data_MPORT_data; // @[SRAM_1.scala 83:25]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_5_en & mem_MPORT_5_mask) begin
      mem[mem_MPORT_5_addr] <= mem_MPORT_5_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_6_en & mem_MPORT_6_mask) begin
      mem[mem_MPORT_6_addr] <= mem_MPORT_6_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_7_en & mem_MPORT_7_mask) begin
      mem[mem_MPORT_7_addr] <= mem_MPORT_7_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_8_en & mem_MPORT_8_mask) begin
      mem[mem_MPORT_8_addr] <= mem_MPORT_8_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_9_en & mem_MPORT_9_mask) begin
      mem[mem_MPORT_9_addr] <= mem_MPORT_9_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_10_en & mem_MPORT_10_mask) begin
      mem[mem_MPORT_10_addr] <= mem_MPORT_10_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_11_en & mem_MPORT_11_mask) begin
      mem[mem_MPORT_11_addr] <= mem_MPORT_11_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_12_en & mem_MPORT_12_mask) begin
      mem[mem_MPORT_12_addr] <= mem_MPORT_12_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_13_en & mem_MPORT_13_mask) begin
      mem[mem_MPORT_13_addr] <= mem_MPORT_13_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_14_en & mem_MPORT_14_mask) begin
      mem[mem_MPORT_14_addr] <= mem_MPORT_14_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_15_en & mem_MPORT_15_mask) begin
      mem[mem_MPORT_15_addr] <= mem_MPORT_15_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_16_en & mem_MPORT_16_mask) begin
      mem[mem_MPORT_16_addr] <= mem_MPORT_16_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_17_en & mem_MPORT_17_mask) begin
      mem[mem_MPORT_17_addr] <= mem_MPORT_17_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_18_en & mem_MPORT_18_mask) begin
      mem[mem_MPORT_18_addr] <= mem_MPORT_18_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_19_en & mem_MPORT_19_mask) begin
      mem[mem_MPORT_19_addr] <= mem_MPORT_19_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_20_en & mem_MPORT_20_mask) begin
      mem[mem_MPORT_20_addr] <= mem_MPORT_20_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_21_en & mem_MPORT_21_mask) begin
      mem[mem_MPORT_21_addr] <= mem_MPORT_21_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_22_en & mem_MPORT_22_mask) begin
      mem[mem_MPORT_22_addr] <= mem_MPORT_22_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_23_en & mem_MPORT_23_mask) begin
      mem[mem_MPORT_23_addr] <= mem_MPORT_23_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_24_en & mem_MPORT_24_mask) begin
      mem[mem_MPORT_24_addr] <= mem_MPORT_24_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_25_en & mem_MPORT_25_mask) begin
      mem[mem_MPORT_25_addr] <= mem_MPORT_25_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_26_en & mem_MPORT_26_mask) begin
      mem[mem_MPORT_26_addr] <= mem_MPORT_26_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_27_en & mem_MPORT_27_mask) begin
      mem[mem_MPORT_27_addr] <= mem_MPORT_27_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_28_en & mem_MPORT_28_mask) begin
      mem[mem_MPORT_28_addr] <= mem_MPORT_28_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_29_en & mem_MPORT_29_mask) begin
      mem[mem_MPORT_29_addr] <= mem_MPORT_29_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_30_en & mem_MPORT_30_mask) begin
      mem[mem_MPORT_30_addr] <= mem_MPORT_30_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_31_en & mem_MPORT_31_mask) begin
      mem[mem_MPORT_31_addr] <= mem_MPORT_31_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_32_en & mem_MPORT_32_mask) begin
      mem[mem_MPORT_32_addr] <= mem_MPORT_32_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_33_en & mem_MPORT_33_mask) begin
      mem[mem_MPORT_33_addr] <= mem_MPORT_33_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_34_en & mem_MPORT_34_mask) begin
      mem[mem_MPORT_34_addr] <= mem_MPORT_34_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_35_en & mem_MPORT_35_mask) begin
      mem[mem_MPORT_35_addr] <= mem_MPORT_35_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_36_en & mem_MPORT_36_mask) begin
      mem[mem_MPORT_36_addr] <= mem_MPORT_36_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_37_en & mem_MPORT_37_mask) begin
      mem[mem_MPORT_37_addr] <= mem_MPORT_37_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_38_en & mem_MPORT_38_mask) begin
      mem[mem_MPORT_38_addr] <= mem_MPORT_38_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_39_en & mem_MPORT_39_mask) begin
      mem[mem_MPORT_39_addr] <= mem_MPORT_39_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_40_en & mem_MPORT_40_mask) begin
      mem[mem_MPORT_40_addr] <= mem_MPORT_40_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_41_en & mem_MPORT_41_mask) begin
      mem[mem_MPORT_41_addr] <= mem_MPORT_41_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_42_en & mem_MPORT_42_mask) begin
      mem[mem_MPORT_42_addr] <= mem_MPORT_42_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_43_en & mem_MPORT_43_mask) begin
      mem[mem_MPORT_43_addr] <= mem_MPORT_43_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_44_en & mem_MPORT_44_mask) begin
      mem[mem_MPORT_44_addr] <= mem_MPORT_44_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_45_en & mem_MPORT_45_mask) begin
      mem[mem_MPORT_45_addr] <= mem_MPORT_45_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_46_en & mem_MPORT_46_mask) begin
      mem[mem_MPORT_46_addr] <= mem_MPORT_46_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_47_en & mem_MPORT_47_mask) begin
      mem[mem_MPORT_47_addr] <= mem_MPORT_47_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_48_en & mem_MPORT_48_mask) begin
      mem[mem_MPORT_48_addr] <= mem_MPORT_48_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_49_en & mem_MPORT_49_mask) begin
      mem[mem_MPORT_49_addr] <= mem_MPORT_49_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_50_en & mem_MPORT_50_mask) begin
      mem[mem_MPORT_50_addr] <= mem_MPORT_50_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_51_en & mem_MPORT_51_mask) begin
      mem[mem_MPORT_51_addr] <= mem_MPORT_51_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_52_en & mem_MPORT_52_mask) begin
      mem[mem_MPORT_52_addr] <= mem_MPORT_52_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_53_en & mem_MPORT_53_mask) begin
      mem[mem_MPORT_53_addr] <= mem_MPORT_53_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_54_en & mem_MPORT_54_mask) begin
      mem[mem_MPORT_54_addr] <= mem_MPORT_54_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_55_en & mem_MPORT_55_mask) begin
      mem[mem_MPORT_55_addr] <= mem_MPORT_55_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_56_en & mem_MPORT_56_mask) begin
      mem[mem_MPORT_56_addr] <= mem_MPORT_56_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_57_en & mem_MPORT_57_mask) begin
      mem[mem_MPORT_57_addr] <= mem_MPORT_57_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_58_en & mem_MPORT_58_mask) begin
      mem[mem_MPORT_58_addr] <= mem_MPORT_58_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_59_en & mem_MPORT_59_mask) begin
      mem[mem_MPORT_59_addr] <= mem_MPORT_59_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_60_en & mem_MPORT_60_mask) begin
      mem[mem_MPORT_60_addr] <= mem_MPORT_60_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_61_en & mem_MPORT_61_mask) begin
      mem[mem_MPORT_61_addr] <= mem_MPORT_61_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_62_en & mem_MPORT_62_mask) begin
      mem[mem_MPORT_62_addr] <= mem_MPORT_62_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_63_en & mem_MPORT_63_mask) begin
      mem[mem_MPORT_63_addr] <= mem_MPORT_63_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_64_en & mem_MPORT_64_mask) begin
      mem[mem_MPORT_64_addr] <= mem_MPORT_64_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_65_en & mem_MPORT_65_mask) begin
      mem[mem_MPORT_65_addr] <= mem_MPORT_65_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_66_en & mem_MPORT_66_mask) begin
      mem[mem_MPORT_66_addr] <= mem_MPORT_66_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_67_en & mem_MPORT_67_mask) begin
      mem[mem_MPORT_67_addr] <= mem_MPORT_67_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_68_en & mem_MPORT_68_mask) begin
      mem[mem_MPORT_68_addr] <= mem_MPORT_68_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_69_en & mem_MPORT_69_mask) begin
      mem[mem_MPORT_69_addr] <= mem_MPORT_69_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_70_en & mem_MPORT_70_mask) begin
      mem[mem_MPORT_70_addr] <= mem_MPORT_70_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_71_en & mem_MPORT_71_mask) begin
      mem[mem_MPORT_71_addr] <= mem_MPORT_71_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_72_en & mem_MPORT_72_mask) begin
      mem[mem_MPORT_72_addr] <= mem_MPORT_72_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_73_en & mem_MPORT_73_mask) begin
      mem[mem_MPORT_73_addr] <= mem_MPORT_73_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_74_en & mem_MPORT_74_mask) begin
      mem[mem_MPORT_74_addr] <= mem_MPORT_74_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_75_en & mem_MPORT_75_mask) begin
      mem[mem_MPORT_75_addr] <= mem_MPORT_75_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_76_en & mem_MPORT_76_mask) begin
      mem[mem_MPORT_76_addr] <= mem_MPORT_76_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_77_en & mem_MPORT_77_mask) begin
      mem[mem_MPORT_77_addr] <= mem_MPORT_77_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_78_en & mem_MPORT_78_mask) begin
      mem[mem_MPORT_78_addr] <= mem_MPORT_78_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_79_en & mem_MPORT_79_mask) begin
      mem[mem_MPORT_79_addr] <= mem_MPORT_79_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_80_en & mem_MPORT_80_mask) begin
      mem[mem_MPORT_80_addr] <= mem_MPORT_80_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_81_en & mem_MPORT_81_mask) begin
      mem[mem_MPORT_81_addr] <= mem_MPORT_81_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_82_en & mem_MPORT_82_mask) begin
      mem[mem_MPORT_82_addr] <= mem_MPORT_82_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_83_en & mem_MPORT_83_mask) begin
      mem[mem_MPORT_83_addr] <= mem_MPORT_83_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_84_en & mem_MPORT_84_mask) begin
      mem[mem_MPORT_84_addr] <= mem_MPORT_84_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_85_en & mem_MPORT_85_mask) begin
      mem[mem_MPORT_85_addr] <= mem_MPORT_85_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_86_en & mem_MPORT_86_mask) begin
      mem[mem_MPORT_86_addr] <= mem_MPORT_86_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_87_en & mem_MPORT_87_mask) begin
      mem[mem_MPORT_87_addr] <= mem_MPORT_87_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_88_en & mem_MPORT_88_mask) begin
      mem[mem_MPORT_88_addr] <= mem_MPORT_88_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_89_en & mem_MPORT_89_mask) begin
      mem[mem_MPORT_89_addr] <= mem_MPORT_89_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_90_en & mem_MPORT_90_mask) begin
      mem[mem_MPORT_90_addr] <= mem_MPORT_90_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_91_en & mem_MPORT_91_mask) begin
      mem[mem_MPORT_91_addr] <= mem_MPORT_91_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_92_en & mem_MPORT_92_mask) begin
      mem[mem_MPORT_92_addr] <= mem_MPORT_92_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_93_en & mem_MPORT_93_mask) begin
      mem[mem_MPORT_93_addr] <= mem_MPORT_93_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_94_en & mem_MPORT_94_mask) begin
      mem[mem_MPORT_94_addr] <= mem_MPORT_94_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_95_en & mem_MPORT_95_mask) begin
      mem[mem_MPORT_95_addr] <= mem_MPORT_95_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_96_en & mem_MPORT_96_mask) begin
      mem[mem_MPORT_96_addr] <= mem_MPORT_96_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_97_en & mem_MPORT_97_mask) begin
      mem[mem_MPORT_97_addr] <= mem_MPORT_97_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_98_en & mem_MPORT_98_mask) begin
      mem[mem_MPORT_98_addr] <= mem_MPORT_98_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_99_en & mem_MPORT_99_mask) begin
      mem[mem_MPORT_99_addr] <= mem_MPORT_99_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_100_en & mem_MPORT_100_mask) begin
      mem[mem_MPORT_100_addr] <= mem_MPORT_100_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_101_en & mem_MPORT_101_mask) begin
      mem[mem_MPORT_101_addr] <= mem_MPORT_101_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_102_en & mem_MPORT_102_mask) begin
      mem[mem_MPORT_102_addr] <= mem_MPORT_102_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_103_en & mem_MPORT_103_mask) begin
      mem[mem_MPORT_103_addr] <= mem_MPORT_103_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_104_en & mem_MPORT_104_mask) begin
      mem[mem_MPORT_104_addr] <= mem_MPORT_104_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_105_en & mem_MPORT_105_mask) begin
      mem[mem_MPORT_105_addr] <= mem_MPORT_105_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_106_en & mem_MPORT_106_mask) begin
      mem[mem_MPORT_106_addr] <= mem_MPORT_106_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_107_en & mem_MPORT_107_mask) begin
      mem[mem_MPORT_107_addr] <= mem_MPORT_107_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_108_en & mem_MPORT_108_mask) begin
      mem[mem_MPORT_108_addr] <= mem_MPORT_108_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_109_en & mem_MPORT_109_mask) begin
      mem[mem_MPORT_109_addr] <= mem_MPORT_109_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_110_en & mem_MPORT_110_mask) begin
      mem[mem_MPORT_110_addr] <= mem_MPORT_110_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_111_en & mem_MPORT_111_mask) begin
      mem[mem_MPORT_111_addr] <= mem_MPORT_111_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_112_en & mem_MPORT_112_mask) begin
      mem[mem_MPORT_112_addr] <= mem_MPORT_112_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_113_en & mem_MPORT_113_mask) begin
      mem[mem_MPORT_113_addr] <= mem_MPORT_113_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_114_en & mem_MPORT_114_mask) begin
      mem[mem_MPORT_114_addr] <= mem_MPORT_114_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_115_en & mem_MPORT_115_mask) begin
      mem[mem_MPORT_115_addr] <= mem_MPORT_115_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_116_en & mem_MPORT_116_mask) begin
      mem[mem_MPORT_116_addr] <= mem_MPORT_116_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_117_en & mem_MPORT_117_mask) begin
      mem[mem_MPORT_117_addr] <= mem_MPORT_117_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_118_en & mem_MPORT_118_mask) begin
      mem[mem_MPORT_118_addr] <= mem_MPORT_118_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_119_en & mem_MPORT_119_mask) begin
      mem[mem_MPORT_119_addr] <= mem_MPORT_119_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_120_en & mem_MPORT_120_mask) begin
      mem[mem_MPORT_120_addr] <= mem_MPORT_120_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_121_en & mem_MPORT_121_mask) begin
      mem[mem_MPORT_121_addr] <= mem_MPORT_121_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_122_en & mem_MPORT_122_mask) begin
      mem[mem_MPORT_122_addr] <= mem_MPORT_122_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_123_en & mem_MPORT_123_mask) begin
      mem[mem_MPORT_123_addr] <= mem_MPORT_123_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_124_en & mem_MPORT_124_mask) begin
      mem[mem_MPORT_124_addr] <= mem_MPORT_124_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_125_en & mem_MPORT_125_mask) begin
      mem[mem_MPORT_125_addr] <= mem_MPORT_125_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_126_en & mem_MPORT_126_mask) begin
      mem[mem_MPORT_126_addr] <= mem_MPORT_126_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_127_en & mem_MPORT_127_mask) begin
      mem[mem_MPORT_127_addr] <= mem_MPORT_127_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_128_en & mem_MPORT_128_mask) begin
      mem[mem_MPORT_128_addr] <= mem_MPORT_128_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_129_en & mem_MPORT_129_mask) begin
      mem[mem_MPORT_129_addr] <= mem_MPORT_129_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_130_en & mem_MPORT_130_mask) begin
      mem[mem_MPORT_130_addr] <= mem_MPORT_130_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_131_en & mem_MPORT_131_mask) begin
      mem[mem_MPORT_131_addr] <= mem_MPORT_131_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_132_en & mem_MPORT_132_mask) begin
      mem[mem_MPORT_132_addr] <= mem_MPORT_132_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_133_en & mem_MPORT_133_mask) begin
      mem[mem_MPORT_133_addr] <= mem_MPORT_133_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_134_en & mem_MPORT_134_mask) begin
      mem[mem_MPORT_134_addr] <= mem_MPORT_134_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_135_en & mem_MPORT_135_mask) begin
      mem[mem_MPORT_135_addr] <= mem_MPORT_135_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_136_en & mem_MPORT_136_mask) begin
      mem[mem_MPORT_136_addr] <= mem_MPORT_136_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_137_en & mem_MPORT_137_mask) begin
      mem[mem_MPORT_137_addr] <= mem_MPORT_137_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_138_en & mem_MPORT_138_mask) begin
      mem[mem_MPORT_138_addr] <= mem_MPORT_138_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_139_en & mem_MPORT_139_mask) begin
      mem[mem_MPORT_139_addr] <= mem_MPORT_139_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_140_en & mem_MPORT_140_mask) begin
      mem[mem_MPORT_140_addr] <= mem_MPORT_140_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_141_en & mem_MPORT_141_mask) begin
      mem[mem_MPORT_141_addr] <= mem_MPORT_141_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_142_en & mem_MPORT_142_mask) begin
      mem[mem_MPORT_142_addr] <= mem_MPORT_142_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_143_en & mem_MPORT_143_mask) begin
      mem[mem_MPORT_143_addr] <= mem_MPORT_143_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_144_en & mem_MPORT_144_mask) begin
      mem[mem_MPORT_144_addr] <= mem_MPORT_144_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_145_en & mem_MPORT_145_mask) begin
      mem[mem_MPORT_145_addr] <= mem_MPORT_145_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_146_en & mem_MPORT_146_mask) begin
      mem[mem_MPORT_146_addr] <= mem_MPORT_146_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_147_en & mem_MPORT_147_mask) begin
      mem[mem_MPORT_147_addr] <= mem_MPORT_147_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_148_en & mem_MPORT_148_mask) begin
      mem[mem_MPORT_148_addr] <= mem_MPORT_148_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_149_en & mem_MPORT_149_mask) begin
      mem[mem_MPORT_149_addr] <= mem_MPORT_149_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_150_en & mem_MPORT_150_mask) begin
      mem[mem_MPORT_150_addr] <= mem_MPORT_150_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_151_en & mem_MPORT_151_mask) begin
      mem[mem_MPORT_151_addr] <= mem_MPORT_151_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_152_en & mem_MPORT_152_mask) begin
      mem[mem_MPORT_152_addr] <= mem_MPORT_152_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_153_en & mem_MPORT_153_mask) begin
      mem[mem_MPORT_153_addr] <= mem_MPORT_153_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_154_en & mem_MPORT_154_mask) begin
      mem[mem_MPORT_154_addr] <= mem_MPORT_154_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_155_en & mem_MPORT_155_mask) begin
      mem[mem_MPORT_155_addr] <= mem_MPORT_155_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_156_en & mem_MPORT_156_mask) begin
      mem[mem_MPORT_156_addr] <= mem_MPORT_156_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_157_en & mem_MPORT_157_mask) begin
      mem[mem_MPORT_157_addr] <= mem_MPORT_157_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_158_en & mem_MPORT_158_mask) begin
      mem[mem_MPORT_158_addr] <= mem_MPORT_158_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_159_en & mem_MPORT_159_mask) begin
      mem[mem_MPORT_159_addr] <= mem_MPORT_159_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_160_en & mem_MPORT_160_mask) begin
      mem[mem_MPORT_160_addr] <= mem_MPORT_160_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_161_en & mem_MPORT_161_mask) begin
      mem[mem_MPORT_161_addr] <= mem_MPORT_161_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_162_en & mem_MPORT_162_mask) begin
      mem[mem_MPORT_162_addr] <= mem_MPORT_162_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_163_en & mem_MPORT_163_mask) begin
      mem[mem_MPORT_163_addr] <= mem_MPORT_163_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_164_en & mem_MPORT_164_mask) begin
      mem[mem_MPORT_164_addr] <= mem_MPORT_164_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_165_en & mem_MPORT_165_mask) begin
      mem[mem_MPORT_165_addr] <= mem_MPORT_165_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_166_en & mem_MPORT_166_mask) begin
      mem[mem_MPORT_166_addr] <= mem_MPORT_166_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_167_en & mem_MPORT_167_mask) begin
      mem[mem_MPORT_167_addr] <= mem_MPORT_167_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_168_en & mem_MPORT_168_mask) begin
      mem[mem_MPORT_168_addr] <= mem_MPORT_168_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_169_en & mem_MPORT_169_mask) begin
      mem[mem_MPORT_169_addr] <= mem_MPORT_169_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_170_en & mem_MPORT_170_mask) begin
      mem[mem_MPORT_170_addr] <= mem_MPORT_170_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_171_en & mem_MPORT_171_mask) begin
      mem[mem_MPORT_171_addr] <= mem_MPORT_171_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_172_en & mem_MPORT_172_mask) begin
      mem[mem_MPORT_172_addr] <= mem_MPORT_172_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_173_en & mem_MPORT_173_mask) begin
      mem[mem_MPORT_173_addr] <= mem_MPORT_173_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_174_en & mem_MPORT_174_mask) begin
      mem[mem_MPORT_174_addr] <= mem_MPORT_174_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_175_en & mem_MPORT_175_mask) begin
      mem[mem_MPORT_175_addr] <= mem_MPORT_175_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_176_en & mem_MPORT_176_mask) begin
      mem[mem_MPORT_176_addr] <= mem_MPORT_176_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_177_en & mem_MPORT_177_mask) begin
      mem[mem_MPORT_177_addr] <= mem_MPORT_177_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_178_en & mem_MPORT_178_mask) begin
      mem[mem_MPORT_178_addr] <= mem_MPORT_178_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_179_en & mem_MPORT_179_mask) begin
      mem[mem_MPORT_179_addr] <= mem_MPORT_179_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_180_en & mem_MPORT_180_mask) begin
      mem[mem_MPORT_180_addr] <= mem_MPORT_180_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_181_en & mem_MPORT_181_mask) begin
      mem[mem_MPORT_181_addr] <= mem_MPORT_181_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_182_en & mem_MPORT_182_mask) begin
      mem[mem_MPORT_182_addr] <= mem_MPORT_182_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_183_en & mem_MPORT_183_mask) begin
      mem[mem_MPORT_183_addr] <= mem_MPORT_183_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_184_en & mem_MPORT_184_mask) begin
      mem[mem_MPORT_184_addr] <= mem_MPORT_184_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_185_en & mem_MPORT_185_mask) begin
      mem[mem_MPORT_185_addr] <= mem_MPORT_185_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_186_en & mem_MPORT_186_mask) begin
      mem[mem_MPORT_186_addr] <= mem_MPORT_186_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_187_en & mem_MPORT_187_mask) begin
      mem[mem_MPORT_187_addr] <= mem_MPORT_187_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_188_en & mem_MPORT_188_mask) begin
      mem[mem_MPORT_188_addr] <= mem_MPORT_188_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_189_en & mem_MPORT_189_mask) begin
      mem[mem_MPORT_189_addr] <= mem_MPORT_189_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_190_en & mem_MPORT_190_mask) begin
      mem[mem_MPORT_190_addr] <= mem_MPORT_190_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_191_en & mem_MPORT_191_mask) begin
      mem[mem_MPORT_191_addr] <= mem_MPORT_191_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_192_en & mem_MPORT_192_mask) begin
      mem[mem_MPORT_192_addr] <= mem_MPORT_192_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_193_en & mem_MPORT_193_mask) begin
      mem[mem_MPORT_193_addr] <= mem_MPORT_193_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_194_en & mem_MPORT_194_mask) begin
      mem[mem_MPORT_194_addr] <= mem_MPORT_194_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_195_en & mem_MPORT_195_mask) begin
      mem[mem_MPORT_195_addr] <= mem_MPORT_195_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_196_en & mem_MPORT_196_mask) begin
      mem[mem_MPORT_196_addr] <= mem_MPORT_196_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_197_en & mem_MPORT_197_mask) begin
      mem[mem_MPORT_197_addr] <= mem_MPORT_197_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_198_en & mem_MPORT_198_mask) begin
      mem[mem_MPORT_198_addr] <= mem_MPORT_198_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_199_en & mem_MPORT_199_mask) begin
      mem[mem_MPORT_199_addr] <= mem_MPORT_199_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_200_en & mem_MPORT_200_mask) begin
      mem[mem_MPORT_200_addr] <= mem_MPORT_200_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_201_en & mem_MPORT_201_mask) begin
      mem[mem_MPORT_201_addr] <= mem_MPORT_201_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_202_en & mem_MPORT_202_mask) begin
      mem[mem_MPORT_202_addr] <= mem_MPORT_202_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_203_en & mem_MPORT_203_mask) begin
      mem[mem_MPORT_203_addr] <= mem_MPORT_203_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_204_en & mem_MPORT_204_mask) begin
      mem[mem_MPORT_204_addr] <= mem_MPORT_204_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_205_en & mem_MPORT_205_mask) begin
      mem[mem_MPORT_205_addr] <= mem_MPORT_205_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_206_en & mem_MPORT_206_mask) begin
      mem[mem_MPORT_206_addr] <= mem_MPORT_206_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_207_en & mem_MPORT_207_mask) begin
      mem[mem_MPORT_207_addr] <= mem_MPORT_207_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_208_en & mem_MPORT_208_mask) begin
      mem[mem_MPORT_208_addr] <= mem_MPORT_208_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_209_en & mem_MPORT_209_mask) begin
      mem[mem_MPORT_209_addr] <= mem_MPORT_209_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_210_en & mem_MPORT_210_mask) begin
      mem[mem_MPORT_210_addr] <= mem_MPORT_210_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_211_en & mem_MPORT_211_mask) begin
      mem[mem_MPORT_211_addr] <= mem_MPORT_211_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_212_en & mem_MPORT_212_mask) begin
      mem[mem_MPORT_212_addr] <= mem_MPORT_212_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_213_en & mem_MPORT_213_mask) begin
      mem[mem_MPORT_213_addr] <= mem_MPORT_213_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_214_en & mem_MPORT_214_mask) begin
      mem[mem_MPORT_214_addr] <= mem_MPORT_214_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_215_en & mem_MPORT_215_mask) begin
      mem[mem_MPORT_215_addr] <= mem_MPORT_215_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_216_en & mem_MPORT_216_mask) begin
      mem[mem_MPORT_216_addr] <= mem_MPORT_216_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_217_en & mem_MPORT_217_mask) begin
      mem[mem_MPORT_217_addr] <= mem_MPORT_217_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_218_en & mem_MPORT_218_mask) begin
      mem[mem_MPORT_218_addr] <= mem_MPORT_218_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_219_en & mem_MPORT_219_mask) begin
      mem[mem_MPORT_219_addr] <= mem_MPORT_219_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_220_en & mem_MPORT_220_mask) begin
      mem[mem_MPORT_220_addr] <= mem_MPORT_220_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_221_en & mem_MPORT_221_mask) begin
      mem[mem_MPORT_221_addr] <= mem_MPORT_221_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_222_en & mem_MPORT_222_mask) begin
      mem[mem_MPORT_222_addr] <= mem_MPORT_222_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_223_en & mem_MPORT_223_mask) begin
      mem[mem_MPORT_223_addr] <= mem_MPORT_223_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_224_en & mem_MPORT_224_mask) begin
      mem[mem_MPORT_224_addr] <= mem_MPORT_224_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_225_en & mem_MPORT_225_mask) begin
      mem[mem_MPORT_225_addr] <= mem_MPORT_225_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_226_en & mem_MPORT_226_mask) begin
      mem[mem_MPORT_226_addr] <= mem_MPORT_226_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_227_en & mem_MPORT_227_mask) begin
      mem[mem_MPORT_227_addr] <= mem_MPORT_227_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_228_en & mem_MPORT_228_mask) begin
      mem[mem_MPORT_228_addr] <= mem_MPORT_228_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_229_en & mem_MPORT_229_mask) begin
      mem[mem_MPORT_229_addr] <= mem_MPORT_229_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_230_en & mem_MPORT_230_mask) begin
      mem[mem_MPORT_230_addr] <= mem_MPORT_230_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_231_en & mem_MPORT_231_mask) begin
      mem[mem_MPORT_231_addr] <= mem_MPORT_231_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_232_en & mem_MPORT_232_mask) begin
      mem[mem_MPORT_232_addr] <= mem_MPORT_232_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_233_en & mem_MPORT_233_mask) begin
      mem[mem_MPORT_233_addr] <= mem_MPORT_233_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_234_en & mem_MPORT_234_mask) begin
      mem[mem_MPORT_234_addr] <= mem_MPORT_234_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_235_en & mem_MPORT_235_mask) begin
      mem[mem_MPORT_235_addr] <= mem_MPORT_235_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_236_en & mem_MPORT_236_mask) begin
      mem[mem_MPORT_236_addr] <= mem_MPORT_236_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_237_en & mem_MPORT_237_mask) begin
      mem[mem_MPORT_237_addr] <= mem_MPORT_237_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_238_en & mem_MPORT_238_mask) begin
      mem[mem_MPORT_238_addr] <= mem_MPORT_238_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_239_en & mem_MPORT_239_mask) begin
      mem[mem_MPORT_239_addr] <= mem_MPORT_239_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_240_en & mem_MPORT_240_mask) begin
      mem[mem_MPORT_240_addr] <= mem_MPORT_240_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_241_en & mem_MPORT_241_mask) begin
      mem[mem_MPORT_241_addr] <= mem_MPORT_241_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_242_en & mem_MPORT_242_mask) begin
      mem[mem_MPORT_242_addr] <= mem_MPORT_242_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_243_en & mem_MPORT_243_mask) begin
      mem[mem_MPORT_243_addr] <= mem_MPORT_243_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_244_en & mem_MPORT_244_mask) begin
      mem[mem_MPORT_244_addr] <= mem_MPORT_244_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_245_en & mem_MPORT_245_mask) begin
      mem[mem_MPORT_245_addr] <= mem_MPORT_245_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_246_en & mem_MPORT_246_mask) begin
      mem[mem_MPORT_246_addr] <= mem_MPORT_246_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_247_en & mem_MPORT_247_mask) begin
      mem[mem_MPORT_247_addr] <= mem_MPORT_247_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_248_en & mem_MPORT_248_mask) begin
      mem[mem_MPORT_248_addr] <= mem_MPORT_248_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_249_en & mem_MPORT_249_mask) begin
      mem[mem_MPORT_249_addr] <= mem_MPORT_249_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_250_en & mem_MPORT_250_mask) begin
      mem[mem_MPORT_250_addr] <= mem_MPORT_250_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_251_en & mem_MPORT_251_mask) begin
      mem[mem_MPORT_251_addr] <= mem_MPORT_251_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_252_en & mem_MPORT_252_mask) begin
      mem[mem_MPORT_252_addr] <= mem_MPORT_252_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_253_en & mem_MPORT_253_mask) begin
      mem[mem_MPORT_253_addr] <= mem_MPORT_253_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_254_en & mem_MPORT_254_mask) begin
      mem[mem_MPORT_254_addr] <= mem_MPORT_254_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_255_en & mem_MPORT_255_mask) begin
      mem[mem_MPORT_255_addr] <= mem_MPORT_255_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_256_en & mem_MPORT_256_mask) begin
      mem[mem_MPORT_256_addr] <= mem_MPORT_256_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_257_en & mem_MPORT_257_mask) begin
      mem[mem_MPORT_257_addr] <= mem_MPORT_257_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_258_en & mem_MPORT_258_mask) begin
      mem[mem_MPORT_258_addr] <= mem_MPORT_258_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_259_en & mem_MPORT_259_mask) begin
      mem[mem_MPORT_259_addr] <= mem_MPORT_259_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_260_en & mem_MPORT_260_mask) begin
      mem[mem_MPORT_260_addr] <= mem_MPORT_260_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_261_en & mem_MPORT_261_mask) begin
      mem[mem_MPORT_261_addr] <= mem_MPORT_261_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_262_en & mem_MPORT_262_mask) begin
      mem[mem_MPORT_262_addr] <= mem_MPORT_262_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_263_en & mem_MPORT_263_mask) begin
      mem[mem_MPORT_263_addr] <= mem_MPORT_263_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_264_en & mem_MPORT_264_mask) begin
      mem[mem_MPORT_264_addr] <= mem_MPORT_264_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_265_en & mem_MPORT_265_mask) begin
      mem[mem_MPORT_265_addr] <= mem_MPORT_265_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_266_en & mem_MPORT_266_mask) begin
      mem[mem_MPORT_266_addr] <= mem_MPORT_266_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_267_en & mem_MPORT_267_mask) begin
      mem[mem_MPORT_267_addr] <= mem_MPORT_267_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_268_en & mem_MPORT_268_mask) begin
      mem[mem_MPORT_268_addr] <= mem_MPORT_268_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_269_en & mem_MPORT_269_mask) begin
      mem[mem_MPORT_269_addr] <= mem_MPORT_269_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_270_en & mem_MPORT_270_mask) begin
      mem[mem_MPORT_270_addr] <= mem_MPORT_270_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_271_en & mem_MPORT_271_mask) begin
      mem[mem_MPORT_271_addr] <= mem_MPORT_271_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_272_en & mem_MPORT_272_mask) begin
      mem[mem_MPORT_272_addr] <= mem_MPORT_272_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_273_en & mem_MPORT_273_mask) begin
      mem[mem_MPORT_273_addr] <= mem_MPORT_273_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_274_en & mem_MPORT_274_mask) begin
      mem[mem_MPORT_274_addr] <= mem_MPORT_274_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_275_en & mem_MPORT_275_mask) begin
      mem[mem_MPORT_275_addr] <= mem_MPORT_275_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_276_en & mem_MPORT_276_mask) begin
      mem[mem_MPORT_276_addr] <= mem_MPORT_276_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_277_en & mem_MPORT_277_mask) begin
      mem[mem_MPORT_277_addr] <= mem_MPORT_277_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_278_en & mem_MPORT_278_mask) begin
      mem[mem_MPORT_278_addr] <= mem_MPORT_278_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_279_en & mem_MPORT_279_mask) begin
      mem[mem_MPORT_279_addr] <= mem_MPORT_279_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_280_en & mem_MPORT_280_mask) begin
      mem[mem_MPORT_280_addr] <= mem_MPORT_280_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_281_en & mem_MPORT_281_mask) begin
      mem[mem_MPORT_281_addr] <= mem_MPORT_281_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_282_en & mem_MPORT_282_mask) begin
      mem[mem_MPORT_282_addr] <= mem_MPORT_282_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_283_en & mem_MPORT_283_mask) begin
      mem[mem_MPORT_283_addr] <= mem_MPORT_283_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_284_en & mem_MPORT_284_mask) begin
      mem[mem_MPORT_284_addr] <= mem_MPORT_284_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_285_en & mem_MPORT_285_mask) begin
      mem[mem_MPORT_285_addr] <= mem_MPORT_285_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_286_en & mem_MPORT_286_mask) begin
      mem[mem_MPORT_286_addr] <= mem_MPORT_286_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_287_en & mem_MPORT_287_mask) begin
      mem[mem_MPORT_287_addr] <= mem_MPORT_287_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_288_en & mem_MPORT_288_mask) begin
      mem[mem_MPORT_288_addr] <= mem_MPORT_288_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_289_en & mem_MPORT_289_mask) begin
      mem[mem_MPORT_289_addr] <= mem_MPORT_289_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_290_en & mem_MPORT_290_mask) begin
      mem[mem_MPORT_290_addr] <= mem_MPORT_290_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_291_en & mem_MPORT_291_mask) begin
      mem[mem_MPORT_291_addr] <= mem_MPORT_291_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_292_en & mem_MPORT_292_mask) begin
      mem[mem_MPORT_292_addr] <= mem_MPORT_292_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_293_en & mem_MPORT_293_mask) begin
      mem[mem_MPORT_293_addr] <= mem_MPORT_293_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_294_en & mem_MPORT_294_mask) begin
      mem[mem_MPORT_294_addr] <= mem_MPORT_294_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_295_en & mem_MPORT_295_mask) begin
      mem[mem_MPORT_295_addr] <= mem_MPORT_295_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_296_en & mem_MPORT_296_mask) begin
      mem[mem_MPORT_296_addr] <= mem_MPORT_296_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_297_en & mem_MPORT_297_mask) begin
      mem[mem_MPORT_297_addr] <= mem_MPORT_297_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_298_en & mem_MPORT_298_mask) begin
      mem[mem_MPORT_298_addr] <= mem_MPORT_298_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_299_en & mem_MPORT_299_mask) begin
      mem[mem_MPORT_299_addr] <= mem_MPORT_299_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_300_en & mem_MPORT_300_mask) begin
      mem[mem_MPORT_300_addr] <= mem_MPORT_300_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_301_en & mem_MPORT_301_mask) begin
      mem[mem_MPORT_301_addr] <= mem_MPORT_301_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_302_en & mem_MPORT_302_mask) begin
      mem[mem_MPORT_302_addr] <= mem_MPORT_302_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_303_en & mem_MPORT_303_mask) begin
      mem[mem_MPORT_303_addr] <= mem_MPORT_303_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_304_en & mem_MPORT_304_mask) begin
      mem[mem_MPORT_304_addr] <= mem_MPORT_304_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_305_en & mem_MPORT_305_mask) begin
      mem[mem_MPORT_305_addr] <= mem_MPORT_305_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_306_en & mem_MPORT_306_mask) begin
      mem[mem_MPORT_306_addr] <= mem_MPORT_306_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_307_en & mem_MPORT_307_mask) begin
      mem[mem_MPORT_307_addr] <= mem_MPORT_307_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_308_en & mem_MPORT_308_mask) begin
      mem[mem_MPORT_308_addr] <= mem_MPORT_308_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_309_en & mem_MPORT_309_mask) begin
      mem[mem_MPORT_309_addr] <= mem_MPORT_309_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_310_en & mem_MPORT_310_mask) begin
      mem[mem_MPORT_310_addr] <= mem_MPORT_310_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_311_en & mem_MPORT_311_mask) begin
      mem[mem_MPORT_311_addr] <= mem_MPORT_311_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_312_en & mem_MPORT_312_mask) begin
      mem[mem_MPORT_312_addr] <= mem_MPORT_312_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_313_en & mem_MPORT_313_mask) begin
      mem[mem_MPORT_313_addr] <= mem_MPORT_313_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_314_en & mem_MPORT_314_mask) begin
      mem[mem_MPORT_314_addr] <= mem_MPORT_314_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_315_en & mem_MPORT_315_mask) begin
      mem[mem_MPORT_315_addr] <= mem_MPORT_315_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_316_en & mem_MPORT_316_mask) begin
      mem[mem_MPORT_316_addr] <= mem_MPORT_316_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_317_en & mem_MPORT_317_mask) begin
      mem[mem_MPORT_317_addr] <= mem_MPORT_317_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_318_en & mem_MPORT_318_mask) begin
      mem[mem_MPORT_318_addr] <= mem_MPORT_318_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_319_en & mem_MPORT_319_mask) begin
      mem[mem_MPORT_319_addr] <= mem_MPORT_319_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_320_en & mem_MPORT_320_mask) begin
      mem[mem_MPORT_320_addr] <= mem_MPORT_320_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_321_en & mem_MPORT_321_mask) begin
      mem[mem_MPORT_321_addr] <= mem_MPORT_321_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_322_en & mem_MPORT_322_mask) begin
      mem[mem_MPORT_322_addr] <= mem_MPORT_322_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_323_en & mem_MPORT_323_mask) begin
      mem[mem_MPORT_323_addr] <= mem_MPORT_323_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_324_en & mem_MPORT_324_mask) begin
      mem[mem_MPORT_324_addr] <= mem_MPORT_324_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_325_en & mem_MPORT_325_mask) begin
      mem[mem_MPORT_325_addr] <= mem_MPORT_325_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_326_en & mem_MPORT_326_mask) begin
      mem[mem_MPORT_326_addr] <= mem_MPORT_326_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_327_en & mem_MPORT_327_mask) begin
      mem[mem_MPORT_327_addr] <= mem_MPORT_327_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_328_en & mem_MPORT_328_mask) begin
      mem[mem_MPORT_328_addr] <= mem_MPORT_328_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_329_en & mem_MPORT_329_mask) begin
      mem[mem_MPORT_329_addr] <= mem_MPORT_329_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_330_en & mem_MPORT_330_mask) begin
      mem[mem_MPORT_330_addr] <= mem_MPORT_330_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_331_en & mem_MPORT_331_mask) begin
      mem[mem_MPORT_331_addr] <= mem_MPORT_331_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_332_en & mem_MPORT_332_mask) begin
      mem[mem_MPORT_332_addr] <= mem_MPORT_332_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_333_en & mem_MPORT_333_mask) begin
      mem[mem_MPORT_333_addr] <= mem_MPORT_333_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_334_en & mem_MPORT_334_mask) begin
      mem[mem_MPORT_334_addr] <= mem_MPORT_334_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_335_en & mem_MPORT_335_mask) begin
      mem[mem_MPORT_335_addr] <= mem_MPORT_335_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_336_en & mem_MPORT_336_mask) begin
      mem[mem_MPORT_336_addr] <= mem_MPORT_336_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_337_en & mem_MPORT_337_mask) begin
      mem[mem_MPORT_337_addr] <= mem_MPORT_337_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_338_en & mem_MPORT_338_mask) begin
      mem[mem_MPORT_338_addr] <= mem_MPORT_338_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_339_en & mem_MPORT_339_mask) begin
      mem[mem_MPORT_339_addr] <= mem_MPORT_339_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_340_en & mem_MPORT_340_mask) begin
      mem[mem_MPORT_340_addr] <= mem_MPORT_340_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_341_en & mem_MPORT_341_mask) begin
      mem[mem_MPORT_341_addr] <= mem_MPORT_341_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_342_en & mem_MPORT_342_mask) begin
      mem[mem_MPORT_342_addr] <= mem_MPORT_342_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_343_en & mem_MPORT_343_mask) begin
      mem[mem_MPORT_343_addr] <= mem_MPORT_343_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_344_en & mem_MPORT_344_mask) begin
      mem[mem_MPORT_344_addr] <= mem_MPORT_344_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_345_en & mem_MPORT_345_mask) begin
      mem[mem_MPORT_345_addr] <= mem_MPORT_345_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_346_en & mem_MPORT_346_mask) begin
      mem[mem_MPORT_346_addr] <= mem_MPORT_346_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_347_en & mem_MPORT_347_mask) begin
      mem[mem_MPORT_347_addr] <= mem_MPORT_347_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_348_en & mem_MPORT_348_mask) begin
      mem[mem_MPORT_348_addr] <= mem_MPORT_348_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_349_en & mem_MPORT_349_mask) begin
      mem[mem_MPORT_349_addr] <= mem_MPORT_349_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_350_en & mem_MPORT_350_mask) begin
      mem[mem_MPORT_350_addr] <= mem_MPORT_350_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_351_en & mem_MPORT_351_mask) begin
      mem[mem_MPORT_351_addr] <= mem_MPORT_351_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_352_en & mem_MPORT_352_mask) begin
      mem[mem_MPORT_352_addr] <= mem_MPORT_352_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_353_en & mem_MPORT_353_mask) begin
      mem[mem_MPORT_353_addr] <= mem_MPORT_353_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_354_en & mem_MPORT_354_mask) begin
      mem[mem_MPORT_354_addr] <= mem_MPORT_354_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_355_en & mem_MPORT_355_mask) begin
      mem[mem_MPORT_355_addr] <= mem_MPORT_355_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_356_en & mem_MPORT_356_mask) begin
      mem[mem_MPORT_356_addr] <= mem_MPORT_356_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_357_en & mem_MPORT_357_mask) begin
      mem[mem_MPORT_357_addr] <= mem_MPORT_357_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_358_en & mem_MPORT_358_mask) begin
      mem[mem_MPORT_358_addr] <= mem_MPORT_358_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_359_en & mem_MPORT_359_mask) begin
      mem[mem_MPORT_359_addr] <= mem_MPORT_359_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_360_en & mem_MPORT_360_mask) begin
      mem[mem_MPORT_360_addr] <= mem_MPORT_360_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_361_en & mem_MPORT_361_mask) begin
      mem[mem_MPORT_361_addr] <= mem_MPORT_361_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_362_en & mem_MPORT_362_mask) begin
      mem[mem_MPORT_362_addr] <= mem_MPORT_362_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_363_en & mem_MPORT_363_mask) begin
      mem[mem_MPORT_363_addr] <= mem_MPORT_363_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_364_en & mem_MPORT_364_mask) begin
      mem[mem_MPORT_364_addr] <= mem_MPORT_364_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_365_en & mem_MPORT_365_mask) begin
      mem[mem_MPORT_365_addr] <= mem_MPORT_365_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_366_en & mem_MPORT_366_mask) begin
      mem[mem_MPORT_366_addr] <= mem_MPORT_366_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_367_en & mem_MPORT_367_mask) begin
      mem[mem_MPORT_367_addr] <= mem_MPORT_367_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_368_en & mem_MPORT_368_mask) begin
      mem[mem_MPORT_368_addr] <= mem_MPORT_368_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_369_en & mem_MPORT_369_mask) begin
      mem[mem_MPORT_369_addr] <= mem_MPORT_369_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_370_en & mem_MPORT_370_mask) begin
      mem[mem_MPORT_370_addr] <= mem_MPORT_370_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_371_en & mem_MPORT_371_mask) begin
      mem[mem_MPORT_371_addr] <= mem_MPORT_371_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_372_en & mem_MPORT_372_mask) begin
      mem[mem_MPORT_372_addr] <= mem_MPORT_372_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_373_en & mem_MPORT_373_mask) begin
      mem[mem_MPORT_373_addr] <= mem_MPORT_373_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_374_en & mem_MPORT_374_mask) begin
      mem[mem_MPORT_374_addr] <= mem_MPORT_374_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_375_en & mem_MPORT_375_mask) begin
      mem[mem_MPORT_375_addr] <= mem_MPORT_375_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_376_en & mem_MPORT_376_mask) begin
      mem[mem_MPORT_376_addr] <= mem_MPORT_376_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_377_en & mem_MPORT_377_mask) begin
      mem[mem_MPORT_377_addr] <= mem_MPORT_377_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_378_en & mem_MPORT_378_mask) begin
      mem[mem_MPORT_378_addr] <= mem_MPORT_378_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_379_en & mem_MPORT_379_mask) begin
      mem[mem_MPORT_379_addr] <= mem_MPORT_379_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_380_en & mem_MPORT_380_mask) begin
      mem[mem_MPORT_380_addr] <= mem_MPORT_380_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_381_en & mem_MPORT_381_mask) begin
      mem[mem_MPORT_381_addr] <= mem_MPORT_381_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_382_en & mem_MPORT_382_mask) begin
      mem[mem_MPORT_382_addr] <= mem_MPORT_382_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_383_en & mem_MPORT_383_mask) begin
      mem[mem_MPORT_383_addr] <= mem_MPORT_383_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_384_en & mem_MPORT_384_mask) begin
      mem[mem_MPORT_384_addr] <= mem_MPORT_384_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_385_en & mem_MPORT_385_mask) begin
      mem[mem_MPORT_385_addr] <= mem_MPORT_385_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_386_en & mem_MPORT_386_mask) begin
      mem[mem_MPORT_386_addr] <= mem_MPORT_386_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_387_en & mem_MPORT_387_mask) begin
      mem[mem_MPORT_387_addr] <= mem_MPORT_387_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_388_en & mem_MPORT_388_mask) begin
      mem[mem_MPORT_388_addr] <= mem_MPORT_388_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_389_en & mem_MPORT_389_mask) begin
      mem[mem_MPORT_389_addr] <= mem_MPORT_389_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_390_en & mem_MPORT_390_mask) begin
      mem[mem_MPORT_390_addr] <= mem_MPORT_390_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_391_en & mem_MPORT_391_mask) begin
      mem[mem_MPORT_391_addr] <= mem_MPORT_391_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_392_en & mem_MPORT_392_mask) begin
      mem[mem_MPORT_392_addr] <= mem_MPORT_392_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_393_en & mem_MPORT_393_mask) begin
      mem[mem_MPORT_393_addr] <= mem_MPORT_393_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_394_en & mem_MPORT_394_mask) begin
      mem[mem_MPORT_394_addr] <= mem_MPORT_394_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_395_en & mem_MPORT_395_mask) begin
      mem[mem_MPORT_395_addr] <= mem_MPORT_395_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_396_en & mem_MPORT_396_mask) begin
      mem[mem_MPORT_396_addr] <= mem_MPORT_396_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_397_en & mem_MPORT_397_mask) begin
      mem[mem_MPORT_397_addr] <= mem_MPORT_397_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_398_en & mem_MPORT_398_mask) begin
      mem[mem_MPORT_398_addr] <= mem_MPORT_398_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_399_en & mem_MPORT_399_mask) begin
      mem[mem_MPORT_399_addr] <= mem_MPORT_399_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_400_en & mem_MPORT_400_mask) begin
      mem[mem_MPORT_400_addr] <= mem_MPORT_400_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_401_en & mem_MPORT_401_mask) begin
      mem[mem_MPORT_401_addr] <= mem_MPORT_401_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_402_en & mem_MPORT_402_mask) begin
      mem[mem_MPORT_402_addr] <= mem_MPORT_402_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_403_en & mem_MPORT_403_mask) begin
      mem[mem_MPORT_403_addr] <= mem_MPORT_403_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_404_en & mem_MPORT_404_mask) begin
      mem[mem_MPORT_404_addr] <= mem_MPORT_404_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_405_en & mem_MPORT_405_mask) begin
      mem[mem_MPORT_405_addr] <= mem_MPORT_405_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_406_en & mem_MPORT_406_mask) begin
      mem[mem_MPORT_406_addr] <= mem_MPORT_406_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_407_en & mem_MPORT_407_mask) begin
      mem[mem_MPORT_407_addr] <= mem_MPORT_407_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_408_en & mem_MPORT_408_mask) begin
      mem[mem_MPORT_408_addr] <= mem_MPORT_408_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_409_en & mem_MPORT_409_mask) begin
      mem[mem_MPORT_409_addr] <= mem_MPORT_409_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_410_en & mem_MPORT_410_mask) begin
      mem[mem_MPORT_410_addr] <= mem_MPORT_410_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_411_en & mem_MPORT_411_mask) begin
      mem[mem_MPORT_411_addr] <= mem_MPORT_411_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_412_en & mem_MPORT_412_mask) begin
      mem[mem_MPORT_412_addr] <= mem_MPORT_412_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_413_en & mem_MPORT_413_mask) begin
      mem[mem_MPORT_413_addr] <= mem_MPORT_413_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_414_en & mem_MPORT_414_mask) begin
      mem[mem_MPORT_414_addr] <= mem_MPORT_414_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_415_en & mem_MPORT_415_mask) begin
      mem[mem_MPORT_415_addr] <= mem_MPORT_415_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_416_en & mem_MPORT_416_mask) begin
      mem[mem_MPORT_416_addr] <= mem_MPORT_416_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_417_en & mem_MPORT_417_mask) begin
      mem[mem_MPORT_417_addr] <= mem_MPORT_417_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_418_en & mem_MPORT_418_mask) begin
      mem[mem_MPORT_418_addr] <= mem_MPORT_418_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_419_en & mem_MPORT_419_mask) begin
      mem[mem_MPORT_419_addr] <= mem_MPORT_419_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_420_en & mem_MPORT_420_mask) begin
      mem[mem_MPORT_420_addr] <= mem_MPORT_420_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_421_en & mem_MPORT_421_mask) begin
      mem[mem_MPORT_421_addr] <= mem_MPORT_421_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_422_en & mem_MPORT_422_mask) begin
      mem[mem_MPORT_422_addr] <= mem_MPORT_422_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_423_en & mem_MPORT_423_mask) begin
      mem[mem_MPORT_423_addr] <= mem_MPORT_423_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_424_en & mem_MPORT_424_mask) begin
      mem[mem_MPORT_424_addr] <= mem_MPORT_424_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_425_en & mem_MPORT_425_mask) begin
      mem[mem_MPORT_425_addr] <= mem_MPORT_425_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_426_en & mem_MPORT_426_mask) begin
      mem[mem_MPORT_426_addr] <= mem_MPORT_426_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_427_en & mem_MPORT_427_mask) begin
      mem[mem_MPORT_427_addr] <= mem_MPORT_427_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_428_en & mem_MPORT_428_mask) begin
      mem[mem_MPORT_428_addr] <= mem_MPORT_428_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_429_en & mem_MPORT_429_mask) begin
      mem[mem_MPORT_429_addr] <= mem_MPORT_429_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_430_en & mem_MPORT_430_mask) begin
      mem[mem_MPORT_430_addr] <= mem_MPORT_430_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_431_en & mem_MPORT_431_mask) begin
      mem[mem_MPORT_431_addr] <= mem_MPORT_431_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_432_en & mem_MPORT_432_mask) begin
      mem[mem_MPORT_432_addr] <= mem_MPORT_432_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_433_en & mem_MPORT_433_mask) begin
      mem[mem_MPORT_433_addr] <= mem_MPORT_433_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_434_en & mem_MPORT_434_mask) begin
      mem[mem_MPORT_434_addr] <= mem_MPORT_434_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_435_en & mem_MPORT_435_mask) begin
      mem[mem_MPORT_435_addr] <= mem_MPORT_435_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_436_en & mem_MPORT_436_mask) begin
      mem[mem_MPORT_436_addr] <= mem_MPORT_436_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_437_en & mem_MPORT_437_mask) begin
      mem[mem_MPORT_437_addr] <= mem_MPORT_437_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_438_en & mem_MPORT_438_mask) begin
      mem[mem_MPORT_438_addr] <= mem_MPORT_438_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_439_en & mem_MPORT_439_mask) begin
      mem[mem_MPORT_439_addr] <= mem_MPORT_439_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_440_en & mem_MPORT_440_mask) begin
      mem[mem_MPORT_440_addr] <= mem_MPORT_440_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_441_en & mem_MPORT_441_mask) begin
      mem[mem_MPORT_441_addr] <= mem_MPORT_441_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_442_en & mem_MPORT_442_mask) begin
      mem[mem_MPORT_442_addr] <= mem_MPORT_442_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_443_en & mem_MPORT_443_mask) begin
      mem[mem_MPORT_443_addr] <= mem_MPORT_443_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_444_en & mem_MPORT_444_mask) begin
      mem[mem_MPORT_444_addr] <= mem_MPORT_444_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_445_en & mem_MPORT_445_mask) begin
      mem[mem_MPORT_445_addr] <= mem_MPORT_445_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_446_en & mem_MPORT_446_mask) begin
      mem[mem_MPORT_446_addr] <= mem_MPORT_446_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_447_en & mem_MPORT_447_mask) begin
      mem[mem_MPORT_447_addr] <= mem_MPORT_447_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_448_en & mem_MPORT_448_mask) begin
      mem[mem_MPORT_448_addr] <= mem_MPORT_448_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_449_en & mem_MPORT_449_mask) begin
      mem[mem_MPORT_449_addr] <= mem_MPORT_449_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_450_en & mem_MPORT_450_mask) begin
      mem[mem_MPORT_450_addr] <= mem_MPORT_450_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_451_en & mem_MPORT_451_mask) begin
      mem[mem_MPORT_451_addr] <= mem_MPORT_451_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_452_en & mem_MPORT_452_mask) begin
      mem[mem_MPORT_452_addr] <= mem_MPORT_452_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_453_en & mem_MPORT_453_mask) begin
      mem[mem_MPORT_453_addr] <= mem_MPORT_453_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_454_en & mem_MPORT_454_mask) begin
      mem[mem_MPORT_454_addr] <= mem_MPORT_454_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_455_en & mem_MPORT_455_mask) begin
      mem[mem_MPORT_455_addr] <= mem_MPORT_455_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_456_en & mem_MPORT_456_mask) begin
      mem[mem_MPORT_456_addr] <= mem_MPORT_456_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_457_en & mem_MPORT_457_mask) begin
      mem[mem_MPORT_457_addr] <= mem_MPORT_457_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_458_en & mem_MPORT_458_mask) begin
      mem[mem_MPORT_458_addr] <= mem_MPORT_458_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_459_en & mem_MPORT_459_mask) begin
      mem[mem_MPORT_459_addr] <= mem_MPORT_459_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_460_en & mem_MPORT_460_mask) begin
      mem[mem_MPORT_460_addr] <= mem_MPORT_460_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_461_en & mem_MPORT_461_mask) begin
      mem[mem_MPORT_461_addr] <= mem_MPORT_461_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_462_en & mem_MPORT_462_mask) begin
      mem[mem_MPORT_462_addr] <= mem_MPORT_462_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_463_en & mem_MPORT_463_mask) begin
      mem[mem_MPORT_463_addr] <= mem_MPORT_463_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_464_en & mem_MPORT_464_mask) begin
      mem[mem_MPORT_464_addr] <= mem_MPORT_464_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_465_en & mem_MPORT_465_mask) begin
      mem[mem_MPORT_465_addr] <= mem_MPORT_465_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_466_en & mem_MPORT_466_mask) begin
      mem[mem_MPORT_466_addr] <= mem_MPORT_466_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_467_en & mem_MPORT_467_mask) begin
      mem[mem_MPORT_467_addr] <= mem_MPORT_467_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_468_en & mem_MPORT_468_mask) begin
      mem[mem_MPORT_468_addr] <= mem_MPORT_468_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_469_en & mem_MPORT_469_mask) begin
      mem[mem_MPORT_469_addr] <= mem_MPORT_469_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_470_en & mem_MPORT_470_mask) begin
      mem[mem_MPORT_470_addr] <= mem_MPORT_470_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_471_en & mem_MPORT_471_mask) begin
      mem[mem_MPORT_471_addr] <= mem_MPORT_471_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_472_en & mem_MPORT_472_mask) begin
      mem[mem_MPORT_472_addr] <= mem_MPORT_472_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_473_en & mem_MPORT_473_mask) begin
      mem[mem_MPORT_473_addr] <= mem_MPORT_473_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_474_en & mem_MPORT_474_mask) begin
      mem[mem_MPORT_474_addr] <= mem_MPORT_474_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_475_en & mem_MPORT_475_mask) begin
      mem[mem_MPORT_475_addr] <= mem_MPORT_475_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_476_en & mem_MPORT_476_mask) begin
      mem[mem_MPORT_476_addr] <= mem_MPORT_476_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_477_en & mem_MPORT_477_mask) begin
      mem[mem_MPORT_477_addr] <= mem_MPORT_477_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_478_en & mem_MPORT_478_mask) begin
      mem[mem_MPORT_478_addr] <= mem_MPORT_478_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_479_en & mem_MPORT_479_mask) begin
      mem[mem_MPORT_479_addr] <= mem_MPORT_479_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_480_en & mem_MPORT_480_mask) begin
      mem[mem_MPORT_480_addr] <= mem_MPORT_480_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_481_en & mem_MPORT_481_mask) begin
      mem[mem_MPORT_481_addr] <= mem_MPORT_481_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_482_en & mem_MPORT_482_mask) begin
      mem[mem_MPORT_482_addr] <= mem_MPORT_482_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_483_en & mem_MPORT_483_mask) begin
      mem[mem_MPORT_483_addr] <= mem_MPORT_483_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_484_en & mem_MPORT_484_mask) begin
      mem[mem_MPORT_484_addr] <= mem_MPORT_484_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_485_en & mem_MPORT_485_mask) begin
      mem[mem_MPORT_485_addr] <= mem_MPORT_485_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_486_en & mem_MPORT_486_mask) begin
      mem[mem_MPORT_486_addr] <= mem_MPORT_486_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_487_en & mem_MPORT_487_mask) begin
      mem[mem_MPORT_487_addr] <= mem_MPORT_487_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_488_en & mem_MPORT_488_mask) begin
      mem[mem_MPORT_488_addr] <= mem_MPORT_488_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_489_en & mem_MPORT_489_mask) begin
      mem[mem_MPORT_489_addr] <= mem_MPORT_489_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_490_en & mem_MPORT_490_mask) begin
      mem[mem_MPORT_490_addr] <= mem_MPORT_490_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_491_en & mem_MPORT_491_mask) begin
      mem[mem_MPORT_491_addr] <= mem_MPORT_491_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_492_en & mem_MPORT_492_mask) begin
      mem[mem_MPORT_492_addr] <= mem_MPORT_492_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_493_en & mem_MPORT_493_mask) begin
      mem[mem_MPORT_493_addr] <= mem_MPORT_493_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_494_en & mem_MPORT_494_mask) begin
      mem[mem_MPORT_494_addr] <= mem_MPORT_494_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_495_en & mem_MPORT_495_mask) begin
      mem[mem_MPORT_495_addr] <= mem_MPORT_495_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_496_en & mem_MPORT_496_mask) begin
      mem[mem_MPORT_496_addr] <= mem_MPORT_496_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_497_en & mem_MPORT_497_mask) begin
      mem[mem_MPORT_497_addr] <= mem_MPORT_497_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_498_en & mem_MPORT_498_mask) begin
      mem[mem_MPORT_498_addr] <= mem_MPORT_498_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_499_en & mem_MPORT_499_mask) begin
      mem[mem_MPORT_499_addr] <= mem_MPORT_499_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_500_en & mem_MPORT_500_mask) begin
      mem[mem_MPORT_500_addr] <= mem_MPORT_500_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_501_en & mem_MPORT_501_mask) begin
      mem[mem_MPORT_501_addr] <= mem_MPORT_501_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_502_en & mem_MPORT_502_mask) begin
      mem[mem_MPORT_502_addr] <= mem_MPORT_502_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_503_en & mem_MPORT_503_mask) begin
      mem[mem_MPORT_503_addr] <= mem_MPORT_503_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_504_en & mem_MPORT_504_mask) begin
      mem[mem_MPORT_504_addr] <= mem_MPORT_504_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_505_en & mem_MPORT_505_mask) begin
      mem[mem_MPORT_505_addr] <= mem_MPORT_505_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_506_en & mem_MPORT_506_mask) begin
      mem[mem_MPORT_506_addr] <= mem_MPORT_506_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_507_en & mem_MPORT_507_mask) begin
      mem[mem_MPORT_507_addr] <= mem_MPORT_507_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_508_en & mem_MPORT_508_mask) begin
      mem[mem_MPORT_508_addr] <= mem_MPORT_508_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_509_en & mem_MPORT_509_mask) begin
      mem[mem_MPORT_509_addr] <= mem_MPORT_509_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_510_en & mem_MPORT_510_mask) begin
      mem[mem_MPORT_510_addr] <= mem_MPORT_510_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_511_en & mem_MPORT_511_mask) begin
      mem[mem_MPORT_511_addr] <= mem_MPORT_511_data; // @[SRAM_1.scala 63:26]
    end
    if (mem_MPORT_512_en & mem_MPORT_512_mask) begin
      mem[mem_MPORT_512_addr] <= mem_MPORT_512_data; // @[SRAM_1.scala 63:26]
    end
    mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
